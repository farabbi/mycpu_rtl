module mul(
  input mul_clk,
  input resetn,
  input mul_signed,
  input [31:0] x,
  input [31:0] y,
  output [63:0] result
);
wire [32:0] x_33bits;
wire [32:0] y_33bits;
assign x_33bits = {x[31] & mul_signed, x};
assign y_33bits = {y[31] & mul_signed, y};

wire [65:0] x_66bits;
assign x_66bits = {{33{x_33bits[32]}}, x_33bits};

wire [65:0] p[16:0];
wire c[16:0];
booth booth_0(
  .x  (x_66bits     ),
  .y0 (1'b0         ),
  .y1 (1'b0         ),
  .y2 (y_33bits[0]  ),
  .p  (p[0]         ),
  .c  (c[0]         )
);
booth booth_1(
  .x  (x_66bits     ),
  .y0 (y_33bits[0]  ),
  .y1 (y_33bits[1]  ),
  .y2 (y_33bits[2]  ),
  .p  (p[1]         ),
  .c  (c[1]         )
);
booth booth_2(
  .x  (x_66bits     ),
  .y0 (y_33bits[2]  ),
  .y1 (y_33bits[3]  ),
  .y2 (y_33bits[4]  ),
  .p  (p[2]         ),
  .c  (c[2]         )
);
booth booth_3(
  .x  (x_66bits     ),
  .y0 (y_33bits[4]  ),
  .y1 (y_33bits[5]  ),
  .y2 (y_33bits[6]  ),
  .p  (p[3]         ),
  .c  (c[3]         )
);
booth booth_4(
  .x  (x_66bits     ),
  .y0 (y_33bits[6]  ),
  .y1 (y_33bits[7]  ),
  .y2 (y_33bits[8]  ),
  .p  (p[4]         ),
  .c  (c[4]         )
);
booth booth_5(
  .x  (x_66bits     ),
  .y0 (y_33bits[8]  ),
  .y1 (y_33bits[9]  ),
  .y2 (y_33bits[10] ),
  .p  (p[5]         ),
  .c  (c[5]         )
);
booth booth_6(
  .x  (x_66bits     ),
  .y0 (y_33bits[10] ),
  .y1 (y_33bits[11] ),
  .y2 (y_33bits[12] ),
  .p  (p[6]         ),
  .c  (c[6]         )
);
booth booth_7(
  .x  (x_66bits     ),
  .y0 (y_33bits[12] ),
  .y1 (y_33bits[13] ),
  .y2 (y_33bits[14] ),
  .p  (p[7]         ),
  .c  (c[7]         )
);
booth booth_8(
  .x  (x_66bits     ),
  .y0 (y_33bits[14] ),
  .y1 (y_33bits[15] ),
  .y2 (y_33bits[16] ),
  .p  (p[8]         ),
  .c  (c[8]         )
);
booth booth_9(
  .x  (x_66bits     ),
  .y0 (y_33bits[16] ),
  .y1 (y_33bits[17] ),
  .y2 (y_33bits[18] ),
  .p  (p[9]         ),
  .c  (c[9]         )
);
booth booth_10(
  .x  (x_66bits     ),
  .y0 (y_33bits[18] ),
  .y1 (y_33bits[19] ),
  .y2 (y_33bits[20] ),
  .p  (p[10]        ),
  .c  (c[10]        )
);
booth booth_11(
  .x  (x_66bits     ),
  .y0 (y_33bits[20] ),
  .y1 (y_33bits[21] ),
  .y2 (y_33bits[22] ),
  .p  (p[11]        ),
  .c  (c[11]        )
);
booth booth_12(
  .x  (x_66bits     ),
  .y0 (y_33bits[22] ),
  .y1 (y_33bits[23] ),
  .y2 (y_33bits[24] ),
  .p  (p[12]        ),
  .c  (c[12]        )
);
booth booth_13(
  .x  (x_66bits     ),
  .y0 (y_33bits[24] ),
  .y1 (y_33bits[25] ),
  .y2 (y_33bits[26] ),
  .p  (p[13]        ),
  .c  (c[13]        )
);
booth booth_14(
  .x  (x_66bits     ),
  .y0 (y_33bits[26] ),
  .y1 (y_33bits[27] ),
  .y2 (y_33bits[28] ),
  .p  (p[14]        ),
  .c  (c[14]        )
);
booth booth_15(
  .x  (x_66bits     ),
  .y0 (y_33bits[28] ),
  .y1 (y_33bits[29] ),
  .y2 (y_33bits[30] ),
  .p  (p[15]        ),
  .c  (c[15]        )
);
booth booth_16(
  .x  (x_66bits     ),
  .y0 (y_33bits[30] ),
  .y1 (y_33bits[31] ),
  .y2 (y_33bits[32] ),
  .p  (p[16]        ),
  .c  (c[16]        )
);

wire [65:0] p_shift[16:0];
wire [16:0] wallace_input[65:0];
assign p_shift[0] = {p[0][65], p[0][65:1]};
assign p_shift[1] = {p[1][64:0], c[1]};
assign p_shift[2] = {p[2][62:0], {3{c[2]}}};
assign p_shift[3] = {p[3][60:0], {5{c[3]}}};
assign p_shift[4] = {p[4][58:0], {7{c[4]}}};
assign p_shift[5] = {p[5][56:0], {9{c[5]}}};
assign p_shift[6] = {p[6][54:0], {11{c[6]}}};
assign p_shift[7] = {p[7][52:0], {13{c[7]}}};
assign p_shift[8] = {p[8][50:0], {15{c[8]}}};
assign p_shift[9] = {p[9][48:0], {17{c[9]}}};
assign p_shift[10] = {p[10][46:0], {19{c[10]}}};
assign p_shift[11] = {p[11][44:0], {21{c[11]}}};
assign p_shift[12] = {p[12][42:0], {23{c[12]}}};
assign p_shift[13] = {p[13][40:0], {25{c[13]}}};
assign p_shift[14] = {p[14][38:0], {27{c[14]}}};
assign p_shift[15] = {p[15][36:0], {29{c[15]}}};
assign p_shift[16] = {p[16][34:0], {31{c[16]}}};
assign wallace_input[0] = {p_shift[0][0], p_shift[1][0], p_shift[2][0],
                           p_shift[3][0], p_shift[4][0], p_shift[5][0],
                           p_shift[6][0], p_shift[7][0], p_shift[8][0],
                           p_shift[9][0], p_shift[10][0], p_shift[11][0],
                           p_shift[12][0], p_shift[13][0], p_shift[14][0],
                           p_shift[15][0], p_shift[16][0]};
assign wallace_input[1] = {p_shift[0][1], p_shift[1][1], p_shift[2][1],
                           p_shift[3][1], p_shift[4][1], p_shift[5][1],
                           p_shift[6][1], p_shift[7][1], p_shift[8][1],
                           p_shift[9][1], p_shift[10][1], p_shift[11][1],
                           p_shift[12][1], p_shift[13][1], p_shift[14][1],
                           p_shift[15][1], p_shift[16][1]};
assign wallace_input[2] = {p_shift[0][2], p_shift[1][2], p_shift[2][2],
                           p_shift[3][2], p_shift[4][2], p_shift[5][2],
                           p_shift[6][2], p_shift[7][2], p_shift[8][2],
                           p_shift[9][2], p_shift[10][2], p_shift[11][2],
                           p_shift[12][2], p_shift[13][2], p_shift[14][2],
                           p_shift[15][2], p_shift[16][2]};
assign wallace_input[3] = {p_shift[0][3], p_shift[1][3], p_shift[2][3],
                           p_shift[3][3], p_shift[4][3], p_shift[5][3],
                           p_shift[6][3], p_shift[7][3], p_shift[8][3],
                           p_shift[9][3], p_shift[10][3], p_shift[11][3],
                           p_shift[12][3], p_shift[13][3], p_shift[14][3],
                           p_shift[15][3], p_shift[16][3]};
assign wallace_input[4] = {p_shift[0][4], p_shift[1][4], p_shift[2][4],
                           p_shift[3][4], p_shift[4][4], p_shift[5][4],
                           p_shift[6][4], p_shift[7][4], p_shift[8][4],
                           p_shift[9][4], p_shift[10][4], p_shift[11][4],
                           p_shift[12][4], p_shift[13][4], p_shift[14][4],
                           p_shift[15][4], p_shift[16][4]};
assign wallace_input[5] = {p_shift[0][5], p_shift[1][5], p_shift[2][5],
                           p_shift[3][5], p_shift[4][5], p_shift[5][5],
                           p_shift[6][5], p_shift[7][5], p_shift[8][5],
                           p_shift[9][5], p_shift[10][5], p_shift[11][5],
                           p_shift[12][5], p_shift[13][5], p_shift[14][5],
                           p_shift[15][5], p_shift[16][5]};
assign wallace_input[6] = {p_shift[0][6], p_shift[1][6], p_shift[2][6],
                           p_shift[3][6], p_shift[4][6], p_shift[5][6],
                           p_shift[6][6], p_shift[7][6], p_shift[8][6],
                           p_shift[9][6], p_shift[10][6], p_shift[11][6],
                           p_shift[12][6], p_shift[13][6], p_shift[14][6],
                           p_shift[15][6], p_shift[16][6]};
assign wallace_input[7] = {p_shift[0][7], p_shift[1][7], p_shift[2][7],
                           p_shift[3][7], p_shift[4][7], p_shift[5][7],
                           p_shift[6][7], p_shift[7][7], p_shift[8][7],
                           p_shift[9][7], p_shift[10][7], p_shift[11][7],
                           p_shift[12][7], p_shift[13][7], p_shift[14][7],
                           p_shift[15][7], p_shift[16][7]};
assign wallace_input[8] = {p_shift[0][8], p_shift[1][8], p_shift[2][8],
                           p_shift[3][8], p_shift[4][8], p_shift[5][8],
                           p_shift[6][8], p_shift[7][8], p_shift[8][8],
                           p_shift[9][8], p_shift[10][8], p_shift[11][8],
                           p_shift[12][8], p_shift[13][8], p_shift[14][8],
                           p_shift[15][8], p_shift[16][8]};
assign wallace_input[9] = {p_shift[0][9], p_shift[1][9], p_shift[2][9],
                           p_shift[3][9], p_shift[4][9], p_shift[5][9],
                           p_shift[6][9], p_shift[7][9], p_shift[8][9],
                           p_shift[9][9], p_shift[10][9], p_shift[11][9],
                           p_shift[12][9], p_shift[13][9], p_shift[14][9],
                           p_shift[15][9], p_shift[16][9]};
assign wallace_input[10] = {p_shift[0][10], p_shift[1][10], p_shift[2][10],
                            p_shift[3][10], p_shift[4][10], p_shift[5][10],
                            p_shift[6][10], p_shift[7][10], p_shift[8][10],
                            p_shift[9][10], p_shift[10][10], p_shift[11][10],
                            p_shift[12][10], p_shift[13][10], p_shift[14][10],
                            p_shift[15][10], p_shift[16][10]};
assign wallace_input[11] = {p_shift[0][11], p_shift[1][11], p_shift[2][11],
                            p_shift[3][11], p_shift[4][11], p_shift[5][11],
                            p_shift[6][11], p_shift[7][11], p_shift[8][11],
                            p_shift[9][11], p_shift[10][11], p_shift[11][11],
                            p_shift[12][11], p_shift[13][11], p_shift[14][11],
                            p_shift[15][11], p_shift[16][11]};
assign wallace_input[12] = {p_shift[0][12], p_shift[1][12], p_shift[2][12],
                            p_shift[3][12], p_shift[4][12], p_shift[5][12],
                            p_shift[6][12], p_shift[7][12], p_shift[8][12],
                            p_shift[9][12], p_shift[10][12], p_shift[11][12],
                            p_shift[12][12], p_shift[13][12], p_shift[14][12],
                            p_shift[15][12], p_shift[16][12]};
assign wallace_input[13] = {p_shift[0][13], p_shift[1][13], p_shift[2][13],
                            p_shift[3][13], p_shift[4][13], p_shift[5][13],
                            p_shift[6][13], p_shift[7][13], p_shift[8][13],
                            p_shift[9][13], p_shift[10][13], p_shift[11][13],
                            p_shift[12][13], p_shift[13][13], p_shift[14][13],
                            p_shift[15][13], p_shift[16][13]};
assign wallace_input[14] = {p_shift[0][14], p_shift[1][14], p_shift[2][14],
                            p_shift[3][14], p_shift[4][14], p_shift[5][14],
                            p_shift[6][14], p_shift[7][14], p_shift[8][14],
                            p_shift[9][14], p_shift[10][14], p_shift[11][14],
                            p_shift[12][14], p_shift[13][14], p_shift[14][14],
                            p_shift[15][14], p_shift[16][14]};
assign wallace_input[15] = {p_shift[0][15], p_shift[1][15], p_shift[2][15],
                            p_shift[3][15], p_shift[4][15], p_shift[5][15],
                            p_shift[6][15], p_shift[7][15], p_shift[8][15],
                            p_shift[9][15], p_shift[10][15], p_shift[11][15],
                            p_shift[12][15], p_shift[13][15], p_shift[14][15],
                            p_shift[15][15], p_shift[16][15]};
assign wallace_input[16] = {p_shift[0][16], p_shift[1][16], p_shift[2][16],
                            p_shift[3][16], p_shift[4][16], p_shift[5][16],
                            p_shift[6][16], p_shift[7][16], p_shift[8][16],
                            p_shift[9][16], p_shift[10][16], p_shift[11][16],
                            p_shift[12][16], p_shift[13][16], p_shift[14][16],
                            p_shift[15][16], p_shift[16][16]};
assign wallace_input[17] = {p_shift[0][17], p_shift[1][17], p_shift[2][17],
                            p_shift[3][17], p_shift[4][17], p_shift[5][17],
                            p_shift[6][17], p_shift[7][17], p_shift[8][17],
                            p_shift[9][17], p_shift[10][17], p_shift[11][17],
                            p_shift[12][17], p_shift[13][17], p_shift[14][17],
                            p_shift[15][17], p_shift[16][17]};
assign wallace_input[18] = {p_shift[0][18], p_shift[1][18], p_shift[2][18],
                            p_shift[3][18], p_shift[4][18], p_shift[5][18],
                            p_shift[6][18], p_shift[7][18], p_shift[8][18],
                            p_shift[9][18], p_shift[10][18], p_shift[11][18],
                            p_shift[12][18], p_shift[13][18], p_shift[14][18],
                            p_shift[15][18], p_shift[16][18]};
assign wallace_input[19] = {p_shift[0][19], p_shift[1][19], p_shift[2][19],
                            p_shift[3][19], p_shift[4][19], p_shift[5][19],
                            p_shift[6][19], p_shift[7][19], p_shift[8][19],
                            p_shift[9][19], p_shift[10][19], p_shift[11][19],
                            p_shift[12][19], p_shift[13][19], p_shift[14][19],
                            p_shift[15][19], p_shift[16][19]};
assign wallace_input[20] = {p_shift[0][20], p_shift[1][20], p_shift[2][20],
                            p_shift[3][20], p_shift[4][20], p_shift[5][20],
                            p_shift[6][20], p_shift[7][20], p_shift[8][20],
                            p_shift[9][20], p_shift[10][20], p_shift[11][20],
                            p_shift[12][20], p_shift[13][20], p_shift[14][20],
                            p_shift[15][20], p_shift[16][20]};
assign wallace_input[21] = {p_shift[0][21], p_shift[1][21], p_shift[2][21],
                            p_shift[3][21], p_shift[4][21], p_shift[5][21],
                            p_shift[6][21], p_shift[7][21], p_shift[8][21],
                            p_shift[9][21], p_shift[10][21], p_shift[11][21],
                            p_shift[12][21], p_shift[13][21], p_shift[14][21],
                            p_shift[15][21], p_shift[16][21]};
assign wallace_input[22] = {p_shift[0][22], p_shift[1][22], p_shift[2][22],
                            p_shift[3][22], p_shift[4][22], p_shift[5][22],
                            p_shift[6][22], p_shift[7][22], p_shift[8][22],
                            p_shift[9][22], p_shift[10][22], p_shift[11][22],
                            p_shift[12][22], p_shift[13][22], p_shift[14][22],
                            p_shift[15][22], p_shift[16][22]};
assign wallace_input[23] = {p_shift[0][23], p_shift[1][23], p_shift[2][23],
                            p_shift[3][23], p_shift[4][23], p_shift[5][23],
                            p_shift[6][23], p_shift[7][23], p_shift[8][23],
                            p_shift[9][23], p_shift[10][23], p_shift[11][23],
                            p_shift[12][23], p_shift[13][23], p_shift[14][23],
                            p_shift[15][23], p_shift[16][23]};
assign wallace_input[24] = {p_shift[0][24], p_shift[1][24], p_shift[2][24],
                            p_shift[3][24], p_shift[4][24], p_shift[5][24],
                            p_shift[6][24], p_shift[7][24], p_shift[8][24],
                            p_shift[9][24], p_shift[10][24], p_shift[11][24],
                            p_shift[12][24], p_shift[13][24], p_shift[14][24],
                            p_shift[15][24], p_shift[16][24]};
assign wallace_input[25] = {p_shift[0][25], p_shift[1][25], p_shift[2][25],
                            p_shift[3][25], p_shift[4][25], p_shift[5][25],
                            p_shift[6][25], p_shift[7][25], p_shift[8][25],
                            p_shift[9][25], p_shift[10][25], p_shift[11][25],
                            p_shift[12][25], p_shift[13][25], p_shift[14][25],
                            p_shift[15][25], p_shift[16][25]};
assign wallace_input[26] = {p_shift[0][26], p_shift[1][26], p_shift[2][26],
                            p_shift[3][26], p_shift[4][26], p_shift[5][26],
                            p_shift[6][26], p_shift[7][26], p_shift[8][26],
                            p_shift[9][26], p_shift[10][26], p_shift[11][26],
                            p_shift[12][26], p_shift[13][26], p_shift[14][26],
                            p_shift[15][26], p_shift[16][26]};
assign wallace_input[27] = {p_shift[0][27], p_shift[1][27], p_shift[2][27],
                            p_shift[3][27], p_shift[4][27], p_shift[5][27],
                            p_shift[6][27], p_shift[7][27], p_shift[8][27],
                            p_shift[9][27], p_shift[10][27], p_shift[11][27],
                            p_shift[12][27], p_shift[13][27], p_shift[14][27],
                            p_shift[15][27], p_shift[16][27]};
assign wallace_input[28] = {p_shift[0][28], p_shift[1][28], p_shift[2][28],
                            p_shift[3][28], p_shift[4][28], p_shift[5][28],
                            p_shift[6][28], p_shift[7][28], p_shift[8][28],
                            p_shift[9][28], p_shift[10][28], p_shift[11][28],
                            p_shift[12][28], p_shift[13][28], p_shift[14][28],
                            p_shift[15][28], p_shift[16][28]};
assign wallace_input[29] = {p_shift[0][29], p_shift[1][29], p_shift[2][29],
                            p_shift[3][29], p_shift[4][29], p_shift[5][29],
                            p_shift[6][29], p_shift[7][29], p_shift[8][29],
                            p_shift[9][29], p_shift[10][29], p_shift[11][29],
                            p_shift[12][29], p_shift[13][29], p_shift[14][29],
                            p_shift[15][29], p_shift[16][29]};
assign wallace_input[30] = {p_shift[0][30], p_shift[1][30], p_shift[2][30],
                            p_shift[3][30], p_shift[4][30], p_shift[5][30],
                            p_shift[6][30], p_shift[7][30], p_shift[8][30],
                            p_shift[9][30], p_shift[10][30], p_shift[11][30],
                            p_shift[12][30], p_shift[13][30], p_shift[14][30],
                            p_shift[15][30], p_shift[16][30]};
assign wallace_input[31] = {p_shift[0][31], p_shift[1][31], p_shift[2][31],
                            p_shift[3][31], p_shift[4][31], p_shift[5][31],
                            p_shift[6][31], p_shift[7][31], p_shift[8][31],
                            p_shift[9][31], p_shift[10][31], p_shift[11][31],
                            p_shift[12][31], p_shift[13][31], p_shift[14][31],
                            p_shift[15][31], p_shift[16][31]};
assign wallace_input[32] = {p_shift[0][32], p_shift[1][32], p_shift[2][32],
                            p_shift[3][32], p_shift[4][32], p_shift[5][32],
                            p_shift[6][32], p_shift[7][32], p_shift[8][32],
                            p_shift[9][32], p_shift[10][32], p_shift[11][32],
                            p_shift[12][32], p_shift[13][32], p_shift[14][32],
                            p_shift[15][32], p_shift[16][32]};
assign wallace_input[33] = {p_shift[0][33], p_shift[1][33], p_shift[2][33],
                            p_shift[3][33], p_shift[4][33], p_shift[5][33],
                            p_shift[6][33], p_shift[7][33], p_shift[8][33],
                            p_shift[9][33], p_shift[10][33], p_shift[11][33],
                            p_shift[12][33], p_shift[13][33], p_shift[14][33],
                            p_shift[15][33], p_shift[16][33]};
assign wallace_input[34] = {p_shift[0][34], p_shift[1][34], p_shift[2][34],
                            p_shift[3][34], p_shift[4][34], p_shift[5][34],
                            p_shift[6][34], p_shift[7][34], p_shift[8][34],
                            p_shift[9][34], p_shift[10][34], p_shift[11][34],
                            p_shift[12][34], p_shift[13][34], p_shift[14][34],
                            p_shift[15][34], p_shift[16][34]};
assign wallace_input[35] = {p_shift[0][35], p_shift[1][35], p_shift[2][35],
                            p_shift[3][35], p_shift[4][35], p_shift[5][35],
                            p_shift[6][35], p_shift[7][35], p_shift[8][35],
                            p_shift[9][35], p_shift[10][35], p_shift[11][35],
                            p_shift[12][35], p_shift[13][35], p_shift[14][35],
                            p_shift[15][35], p_shift[16][35]};
assign wallace_input[36] = {p_shift[0][36], p_shift[1][36], p_shift[2][36],
                            p_shift[3][36], p_shift[4][36], p_shift[5][36],
                            p_shift[6][36], p_shift[7][36], p_shift[8][36],
                            p_shift[9][36], p_shift[10][36], p_shift[11][36],
                            p_shift[12][36], p_shift[13][36], p_shift[14][36],
                            p_shift[15][36], p_shift[16][36]};
assign wallace_input[37] = {p_shift[0][37], p_shift[1][37], p_shift[2][37],
                            p_shift[3][37], p_shift[4][37], p_shift[5][37],
                            p_shift[6][37], p_shift[7][37], p_shift[8][37],
                            p_shift[9][37], p_shift[10][37], p_shift[11][37],
                            p_shift[12][37], p_shift[13][37], p_shift[14][37],
                            p_shift[15][37], p_shift[16][37]};
assign wallace_input[38] = {p_shift[0][38], p_shift[1][38], p_shift[2][38],
                            p_shift[3][38], p_shift[4][38], p_shift[5][38],
                            p_shift[6][38], p_shift[7][38], p_shift[8][38],
                            p_shift[9][38], p_shift[10][38], p_shift[11][38],
                            p_shift[12][38], p_shift[13][38], p_shift[14][38],
                            p_shift[15][38], p_shift[16][38]};
assign wallace_input[39] = {p_shift[0][39], p_shift[1][39], p_shift[2][39],
                            p_shift[3][39], p_shift[4][39], p_shift[5][39],
                            p_shift[6][39], p_shift[7][39], p_shift[8][39],
                            p_shift[9][39], p_shift[10][39], p_shift[11][39],
                            p_shift[12][39], p_shift[13][39], p_shift[14][39],
                            p_shift[15][39], p_shift[16][39]};
assign wallace_input[40] = {p_shift[0][40], p_shift[1][40], p_shift[2][40],
                            p_shift[3][40], p_shift[4][40], p_shift[5][40],
                            p_shift[6][40], p_shift[7][40], p_shift[8][40],
                            p_shift[9][40], p_shift[10][40], p_shift[11][40],
                            p_shift[12][40], p_shift[13][40], p_shift[14][40],
                            p_shift[15][40], p_shift[16][40]};
assign wallace_input[41] = {p_shift[0][41], p_shift[1][41], p_shift[2][41],
                            p_shift[3][41], p_shift[4][41], p_shift[5][41],
                            p_shift[6][41], p_shift[7][41], p_shift[8][41],
                            p_shift[9][41], p_shift[10][41], p_shift[11][41],
                            p_shift[12][41], p_shift[13][41], p_shift[14][41],
                            p_shift[15][41], p_shift[16][41]};
assign wallace_input[42] = {p_shift[0][42], p_shift[1][42], p_shift[2][42],
                            p_shift[3][42], p_shift[4][42], p_shift[5][42],
                            p_shift[6][42], p_shift[7][42], p_shift[8][42],
                            p_shift[9][42], p_shift[10][42], p_shift[11][42],
                            p_shift[12][42], p_shift[13][42], p_shift[14][42],
                            p_shift[15][42], p_shift[16][42]};
assign wallace_input[43] = {p_shift[0][43], p_shift[1][43], p_shift[2][43],
                            p_shift[3][43], p_shift[4][43], p_shift[5][43],
                            p_shift[6][43], p_shift[7][43], p_shift[8][43],
                            p_shift[9][43], p_shift[10][43], p_shift[11][43],
                            p_shift[12][43], p_shift[13][43], p_shift[14][43],
                            p_shift[15][43], p_shift[16][43]};
assign wallace_input[44] = {p_shift[0][44], p_shift[1][44], p_shift[2][44],
                            p_shift[3][44], p_shift[4][44], p_shift[5][44],
                            p_shift[6][44], p_shift[7][44], p_shift[8][44],
                            p_shift[9][44], p_shift[10][44], p_shift[11][44],
                            p_shift[12][44], p_shift[13][44], p_shift[14][44],
                            p_shift[15][44], p_shift[16][44]};
assign wallace_input[45] = {p_shift[0][45], p_shift[1][45], p_shift[2][45],
                            p_shift[3][45], p_shift[4][45], p_shift[5][45],
                            p_shift[6][45], p_shift[7][45], p_shift[8][45],
                            p_shift[9][45], p_shift[10][45], p_shift[11][45],
                            p_shift[12][45], p_shift[13][45], p_shift[14][45],
                            p_shift[15][45], p_shift[16][45]};
assign wallace_input[46] = {p_shift[0][46], p_shift[1][46], p_shift[2][46],
                            p_shift[3][46], p_shift[4][46], p_shift[5][46],
                            p_shift[6][46], p_shift[7][46], p_shift[8][46],
                            p_shift[9][46], p_shift[10][46], p_shift[11][46],
                            p_shift[12][46], p_shift[13][46], p_shift[14][46],
                            p_shift[15][46], p_shift[16][46]};
assign wallace_input[47] = {p_shift[0][47], p_shift[1][47], p_shift[2][47],
                            p_shift[3][47], p_shift[4][47], p_shift[5][47],
                            p_shift[6][47], p_shift[7][47], p_shift[8][47],
                            p_shift[9][47], p_shift[10][47], p_shift[11][47],
                            p_shift[12][47], p_shift[13][47], p_shift[14][47],
                            p_shift[15][47], p_shift[16][47]};
assign wallace_input[48] = {p_shift[0][48], p_shift[1][48], p_shift[2][48],
                            p_shift[3][48], p_shift[4][48], p_shift[5][48],
                            p_shift[6][48], p_shift[7][48], p_shift[8][48],
                            p_shift[9][48], p_shift[10][48], p_shift[11][48],
                            p_shift[12][48], p_shift[13][48], p_shift[14][48],
                            p_shift[15][48], p_shift[16][48]};
assign wallace_input[49] = {p_shift[0][49], p_shift[1][49], p_shift[2][49],
                            p_shift[3][49], p_shift[4][49], p_shift[5][49],
                            p_shift[6][49], p_shift[7][49], p_shift[8][49],
                            p_shift[9][49], p_shift[10][49], p_shift[11][49],
                            p_shift[12][49], p_shift[13][49], p_shift[14][49],
                            p_shift[15][49], p_shift[16][49]};
assign wallace_input[50] = {p_shift[0][50], p_shift[1][50], p_shift[2][50],
                            p_shift[3][50], p_shift[4][50], p_shift[5][50],
                            p_shift[6][50], p_shift[7][50], p_shift[8][50],
                            p_shift[9][50], p_shift[10][50], p_shift[11][50],
                            p_shift[12][50], p_shift[13][50], p_shift[14][50],
                            p_shift[15][50], p_shift[16][50]};
assign wallace_input[51] = {p_shift[0][51], p_shift[1][51], p_shift[2][51],
                            p_shift[3][51], p_shift[4][51], p_shift[5][51],
                            p_shift[6][51], p_shift[7][51], p_shift[8][51],
                            p_shift[9][51], p_shift[10][51], p_shift[11][51],
                            p_shift[12][51], p_shift[13][51], p_shift[14][51],
                            p_shift[15][51], p_shift[16][51]};
assign wallace_input[52] = {p_shift[0][52], p_shift[1][52], p_shift[2][52],
                            p_shift[3][52], p_shift[4][52], p_shift[5][52],
                            p_shift[6][52], p_shift[7][52], p_shift[8][52],
                            p_shift[9][52], p_shift[10][52], p_shift[11][52],
                            p_shift[12][52], p_shift[13][52], p_shift[14][52],
                            p_shift[15][52], p_shift[16][52]};
assign wallace_input[53] = {p_shift[0][53], p_shift[1][53], p_shift[2][53],
                            p_shift[3][53], p_shift[4][53], p_shift[5][53],
                            p_shift[6][53], p_shift[7][53], p_shift[8][53],
                            p_shift[9][53], p_shift[10][53], p_shift[11][53],
                            p_shift[12][53], p_shift[13][53], p_shift[14][53],
                            p_shift[15][53], p_shift[16][53]};
assign wallace_input[54] = {p_shift[0][54], p_shift[1][54], p_shift[2][54],
                            p_shift[3][54], p_shift[4][54], p_shift[5][54],
                            p_shift[6][54], p_shift[7][54], p_shift[8][54],
                            p_shift[9][54], p_shift[10][54], p_shift[11][54],
                            p_shift[12][54], p_shift[13][54], p_shift[14][54],
                            p_shift[15][54], p_shift[16][54]};
assign wallace_input[55] = {p_shift[0][55], p_shift[1][55], p_shift[2][55],
                            p_shift[3][55], p_shift[4][55], p_shift[5][55],
                            p_shift[6][55], p_shift[7][55], p_shift[8][55],
                            p_shift[9][55], p_shift[10][55], p_shift[11][55],
                            p_shift[12][55], p_shift[13][55], p_shift[14][55],
                            p_shift[15][55], p_shift[16][55]};
assign wallace_input[56] = {p_shift[0][56], p_shift[1][56], p_shift[2][56],
                            p_shift[3][56], p_shift[4][56], p_shift[5][56],
                            p_shift[6][56], p_shift[7][56], p_shift[8][56],
                            p_shift[9][56], p_shift[10][56], p_shift[11][56],
                            p_shift[12][56], p_shift[13][56], p_shift[14][56],
                            p_shift[15][56], p_shift[16][56]};
assign wallace_input[57] = {p_shift[0][57], p_shift[1][57], p_shift[2][57],
                            p_shift[3][57], p_shift[4][57], p_shift[5][57],
                            p_shift[6][57], p_shift[7][57], p_shift[8][57],
                            p_shift[9][57], p_shift[10][57], p_shift[11][57],
                            p_shift[12][57], p_shift[13][57], p_shift[14][57],
                            p_shift[15][57], p_shift[16][57]};
assign wallace_input[58] = {p_shift[0][58], p_shift[1][58], p_shift[2][58],
                            p_shift[3][58], p_shift[4][58], p_shift[5][58],
                            p_shift[6][58], p_shift[7][58], p_shift[8][58],
                            p_shift[9][58], p_shift[10][58], p_shift[11][58],
                            p_shift[12][58], p_shift[13][58], p_shift[14][58],
                            p_shift[15][58], p_shift[16][58]};
assign wallace_input[59] = {p_shift[0][59], p_shift[1][59], p_shift[2][59],
                            p_shift[3][59], p_shift[4][59], p_shift[5][59],
                            p_shift[6][59], p_shift[7][59], p_shift[8][59],
                            p_shift[9][59], p_shift[10][59], p_shift[11][59],
                            p_shift[12][59], p_shift[13][59], p_shift[14][59],
                            p_shift[15][59], p_shift[16][59]};
assign wallace_input[60] = {p_shift[0][60], p_shift[1][60], p_shift[2][60],
                            p_shift[3][60], p_shift[4][60], p_shift[5][60],
                            p_shift[6][60], p_shift[7][60], p_shift[8][60],
                            p_shift[9][60], p_shift[10][60], p_shift[11][60],
                            p_shift[12][60], p_shift[13][60], p_shift[14][60],
                            p_shift[15][60], p_shift[16][60]};
assign wallace_input[61] = {p_shift[0][61], p_shift[1][61], p_shift[2][61],
                            p_shift[3][61], p_shift[4][61], p_shift[5][61],
                            p_shift[6][61], p_shift[7][61], p_shift[8][61],
                            p_shift[9][61], p_shift[10][61], p_shift[11][61],
                            p_shift[12][61], p_shift[13][61], p_shift[14][61],
                            p_shift[15][61], p_shift[16][61]};
assign wallace_input[62] = {p_shift[0][62], p_shift[1][62], p_shift[2][62],
                            p_shift[3][62], p_shift[4][62], p_shift[5][62],
                            p_shift[6][62], p_shift[7][62], p_shift[8][62],
                            p_shift[9][62], p_shift[10][62], p_shift[11][62],
                            p_shift[12][62], p_shift[13][62], p_shift[14][62],
                            p_shift[15][62], p_shift[16][62]};
assign wallace_input[63] = {p_shift[0][63], p_shift[1][63], p_shift[2][63],
                            p_shift[3][63], p_shift[4][63], p_shift[5][63],
                            p_shift[6][63], p_shift[7][63], p_shift[8][63],
                            p_shift[9][63], p_shift[10][63], p_shift[11][63],
                            p_shift[12][63], p_shift[13][63], p_shift[14][63],
                            p_shift[15][63], p_shift[16][63]};
assign wallace_input[64] = {p_shift[0][64], p_shift[1][64], p_shift[2][64],
                            p_shift[3][64], p_shift[4][64], p_shift[5][64],
                            p_shift[6][64], p_shift[7][64], p_shift[8][64],
                            p_shift[9][64], p_shift[10][64], p_shift[11][64],
                            p_shift[12][64], p_shift[13][64], p_shift[14][64],
                            p_shift[15][64], p_shift[16][64]};
assign wallace_input[65] = {p_shift[0][65], p_shift[1][65], p_shift[2][65],
                            p_shift[3][65], p_shift[4][65], p_shift[5][65],
                            p_shift[6][65], p_shift[7][65], p_shift[8][65],
                            p_shift[9][65], p_shift[10][65], p_shift[11][65],
                            p_shift[12][65], p_shift[13][65], p_shift[14][65],
                            p_shift[15][65], p_shift[16][65]};

wire wallace_c[64:0];
wire wallace_s[65:0];
wire [14:0] wallace_cout[64:0];
wallace_tree wallace_tree_0(
	.wallace_input	(wallace_input[0]	),
	.cin_0			(c[0]				),
	.cin_1			(c[1]				),
	.cin_2			(c[2]				),
	.cin_3			(c[3]				),
	.cin_4			(c[4]				),
	.cin_5			(c[5]				),
	.cin_6			(c[6]				),
	.cin_7			(c[7]				),
	.cin_8			(c[8]				),
	.cin_9			(c[9]				),
	.cin_10			(c[10]				),
	.cin_11			(c[11]				),
	.cin_12			(c[12]				),
	.cin_13			(c[13]				),
	.cin_14			(c[14]				),
	.cout_0			(wallace_cout[0][0]	),
	.cout_1			(wallace_cout[0][1]	),
	.cout_2			(wallace_cout[0][2]	),
	.cout_3			(wallace_cout[0][3]	),
	.cout_4			(wallace_cout[0][4]	),
	.cout_5			(wallace_cout[0][5]	),
	.cout_6			(wallace_cout[0][6]	),
	.cout_7			(wallace_cout[0][7]	),
	.cout_8			(wallace_cout[0][8]	),
	.cout_9			(wallace_cout[0][9]	),
	.cout_10		(wallace_cout[0][10]),
	.cout_11		(wallace_cout[0][11]),
	.cout_12		(wallace_cout[0][12]),
	.cout_13		(wallace_cout[0][13]),
	.cout_14		(wallace_cout[0][14]),
	.wallace_c		(wallace_c[0]		),
	.wallace_s		(wallace_s[0]		)
);
wallace_tree wallace_tree_1(
	.wallace_input	(wallace_input[1]	),
	.cin_0			(wallace_cout[0][0] ),
	.cin_1			(wallace_cout[0][1] ),
	.cin_2			(wallace_cout[0][2] ),
	.cin_3			(wallace_cout[0][3] ),
	.cin_4			(wallace_cout[0][4] ),
	.cin_5			(wallace_cout[0][5] ),
	.cin_6			(wallace_cout[0][6] ),
	.cin_7			(wallace_cout[0][7] ),
	.cin_8			(wallace_cout[0][8] ),
	.cin_9			(wallace_cout[0][9] ),
	.cin_10			(wallace_cout[0][10]),
	.cin_11			(wallace_cout[0][11]),
	.cin_12			(wallace_cout[0][12]),
	.cin_13			(wallace_cout[0][13]),
	.cin_14			(wallace_cout[0][14]),
	.cout_0			(wallace_cout[1][0] ),
	.cout_1			(wallace_cout[1][1] ),
	.cout_2			(wallace_cout[1][2] ),
	.cout_3			(wallace_cout[1][3] ),
	.cout_4			(wallace_cout[1][4] ),
	.cout_5			(wallace_cout[1][5] ),
	.cout_6			(wallace_cout[1][6] ),
	.cout_7			(wallace_cout[1][7] ),
	.cout_8			(wallace_cout[1][8] ),
	.cout_9			(wallace_cout[1][9] ),
	.cout_10		(wallace_cout[1][10]),
	.cout_11		(wallace_cout[1][11]),
	.cout_12		(wallace_cout[1][12]),
	.cout_13		(wallace_cout[1][13]),
	.cout_14		(wallace_cout[1][14]),
	.wallace_c		(wallace_c[1]		),
	.wallace_s		(wallace_s[1]		)
);
wallace_tree wallace_tree_2(
	.wallace_input	(wallace_input[2]	),
	.cin_0			(wallace_cout[1][0] ),
	.cin_1			(wallace_cout[1][1] ),
	.cin_2			(wallace_cout[1][2] ),
	.cin_3			(wallace_cout[1][3] ),
	.cin_4			(wallace_cout[1][4] ),
	.cin_5			(wallace_cout[1][5] ),
	.cin_6			(wallace_cout[1][6] ),
	.cin_7			(wallace_cout[1][7] ),
	.cin_8			(wallace_cout[1][8] ),
	.cin_9			(wallace_cout[1][9] ),
	.cin_10			(wallace_cout[1][10]),
	.cin_11			(wallace_cout[1][11]),
	.cin_12			(wallace_cout[1][12]),
	.cin_13			(wallace_cout[1][13]),
	.cin_14			(wallace_cout[1][14]),
	.cout_0			(wallace_cout[2][0] ),
	.cout_1			(wallace_cout[2][1] ),
	.cout_2			(wallace_cout[2][2] ),
	.cout_3			(wallace_cout[2][3] ),
	.cout_4			(wallace_cout[2][4] ),
	.cout_5			(wallace_cout[2][5] ),
	.cout_6			(wallace_cout[2][6] ),
	.cout_7			(wallace_cout[2][7] ),
	.cout_8			(wallace_cout[2][8] ),
	.cout_9			(wallace_cout[2][9] ),
	.cout_10		(wallace_cout[2][10]),
	.cout_11		(wallace_cout[2][11]),
	.cout_12		(wallace_cout[2][12]),
	.cout_13		(wallace_cout[2][13]),
	.cout_14		(wallace_cout[2][14]),
	.wallace_c		(wallace_c[2]		),
	.wallace_s		(wallace_s[2]		)
);
wallace_tree wallace_tree_3(
	.wallace_input	(wallace_input[3]	),
	.cin_0			(wallace_cout[2][0] ),
	.cin_1			(wallace_cout[2][1] ),
	.cin_2			(wallace_cout[2][2] ),
	.cin_3			(wallace_cout[2][3] ),
	.cin_4			(wallace_cout[2][4] ),
	.cin_5			(wallace_cout[2][5] ),
	.cin_6			(wallace_cout[2][6] ),
	.cin_7			(wallace_cout[2][7] ),
	.cin_8			(wallace_cout[2][8] ),
	.cin_9			(wallace_cout[2][9] ),
	.cin_10			(wallace_cout[2][10]),
	.cin_11			(wallace_cout[2][11]),
	.cin_12			(wallace_cout[2][12]),
	.cin_13			(wallace_cout[2][13]),
	.cin_14			(wallace_cout[2][14]),
	.cout_0			(wallace_cout[3][0] ),
	.cout_1			(wallace_cout[3][1] ),
	.cout_2			(wallace_cout[3][2] ),
	.cout_3			(wallace_cout[3][3] ),
	.cout_4			(wallace_cout[3][4] ),
	.cout_5			(wallace_cout[3][5] ),
	.cout_6			(wallace_cout[3][6] ),
	.cout_7			(wallace_cout[3][7] ),
	.cout_8			(wallace_cout[3][8] ),
	.cout_9			(wallace_cout[3][9] ),
	.cout_10		(wallace_cout[3][10]),
	.cout_11		(wallace_cout[3][11]),
	.cout_12		(wallace_cout[3][12]),
	.cout_13		(wallace_cout[3][13]),
	.cout_14		(wallace_cout[3][14]),
	.wallace_c		(wallace_c[3]		),
	.wallace_s		(wallace_s[3]		)
);
wallace_tree wallace_tree_4(
	.wallace_input	(wallace_input[4]	),
	.cin_0			(wallace_cout[3][0] ),
	.cin_1			(wallace_cout[3][1] ),
	.cin_2			(wallace_cout[3][2] ),
	.cin_3			(wallace_cout[3][3] ),
	.cin_4			(wallace_cout[3][4] ),
	.cin_5			(wallace_cout[3][5] ),
	.cin_6			(wallace_cout[3][6] ),
	.cin_7			(wallace_cout[3][7] ),
	.cin_8			(wallace_cout[3][8] ),
	.cin_9			(wallace_cout[3][9] ),
	.cin_10			(wallace_cout[3][10]),
	.cin_11			(wallace_cout[3][11]),
	.cin_12			(wallace_cout[3][12]),
	.cin_13			(wallace_cout[3][13]),
	.cin_14			(wallace_cout[3][14]),
	.cout_0			(wallace_cout[4][0] ),
	.cout_1			(wallace_cout[4][1] ),
	.cout_2			(wallace_cout[4][2] ),
	.cout_3			(wallace_cout[4][3] ),
	.cout_4			(wallace_cout[4][4] ),
	.cout_5			(wallace_cout[4][5] ),
	.cout_6			(wallace_cout[4][6] ),
	.cout_7			(wallace_cout[4][7] ),
	.cout_8			(wallace_cout[4][8] ),
	.cout_9			(wallace_cout[4][9] ),
	.cout_10		(wallace_cout[4][10]),
	.cout_11		(wallace_cout[4][11]),
	.cout_12		(wallace_cout[4][12]),
	.cout_13		(wallace_cout[4][13]),
	.cout_14		(wallace_cout[4][14]),
	.wallace_c		(wallace_c[4]		),
	.wallace_s		(wallace_s[4]		)
);
wallace_tree wallace_tree_5(
	.wallace_input	(wallace_input[5]	),
	.cin_0			(wallace_cout[4][0] ),
	.cin_1			(wallace_cout[4][1] ),
	.cin_2			(wallace_cout[4][2] ),
	.cin_3			(wallace_cout[4][3] ),
	.cin_4			(wallace_cout[4][4] ),
	.cin_5			(wallace_cout[4][5] ),
	.cin_6			(wallace_cout[4][6] ),
	.cin_7			(wallace_cout[4][7] ),
	.cin_8			(wallace_cout[4][8] ),
	.cin_9			(wallace_cout[4][9] ),
	.cin_10			(wallace_cout[4][10]),
	.cin_11			(wallace_cout[4][11]),
	.cin_12			(wallace_cout[4][12]),
	.cin_13			(wallace_cout[4][13]),
	.cin_14			(wallace_cout[4][14]),
	.cout_0			(wallace_cout[5][0] ),
	.cout_1			(wallace_cout[5][1] ),
	.cout_2			(wallace_cout[5][2] ),
	.cout_3			(wallace_cout[5][3] ),
	.cout_4			(wallace_cout[5][4] ),
	.cout_5			(wallace_cout[5][5] ),
	.cout_6			(wallace_cout[5][6] ),
	.cout_7			(wallace_cout[5][7] ),
	.cout_8			(wallace_cout[5][8] ),
	.cout_9			(wallace_cout[5][9] ),
	.cout_10		(wallace_cout[5][10]),
	.cout_11		(wallace_cout[5][11]),
	.cout_12		(wallace_cout[5][12]),
	.cout_13		(wallace_cout[5][13]),
	.cout_14		(wallace_cout[5][14]),
	.wallace_c		(wallace_c[5]		),
	.wallace_s		(wallace_s[5]		)
);
wallace_tree wallace_tree_6(
	.wallace_input	(wallace_input[6]	),
	.cin_0			(wallace_cout[5][0] ),
	.cin_1			(wallace_cout[5][1] ),
	.cin_2			(wallace_cout[5][2] ),
	.cin_3			(wallace_cout[5][3] ),
	.cin_4			(wallace_cout[5][4] ),
	.cin_5			(wallace_cout[5][5] ),
	.cin_6			(wallace_cout[5][6] ),
	.cin_7			(wallace_cout[5][7] ),
	.cin_8			(wallace_cout[5][8] ),
	.cin_9			(wallace_cout[5][9] ),
	.cin_10			(wallace_cout[5][10]),
	.cin_11			(wallace_cout[5][11]),
	.cin_12			(wallace_cout[5][12]),
	.cin_13			(wallace_cout[5][13]),
	.cin_14			(wallace_cout[5][14]),
	.cout_0			(wallace_cout[6][0] ),
	.cout_1			(wallace_cout[6][1] ),
	.cout_2			(wallace_cout[6][2] ),
	.cout_3			(wallace_cout[6][3] ),
	.cout_4			(wallace_cout[6][4] ),
	.cout_5			(wallace_cout[6][5] ),
	.cout_6			(wallace_cout[6][6] ),
	.cout_7			(wallace_cout[6][7] ),
	.cout_8			(wallace_cout[6][8] ),
	.cout_9			(wallace_cout[6][9] ),
	.cout_10		(wallace_cout[6][10]),
	.cout_11		(wallace_cout[6][11]),
	.cout_12		(wallace_cout[6][12]),
	.cout_13		(wallace_cout[6][13]),
	.cout_14		(wallace_cout[6][14]),
	.wallace_c		(wallace_c[6]		),
	.wallace_s		(wallace_s[6]		)
);
wallace_tree wallace_tree_7(
	.wallace_input	(wallace_input[7]	),
	.cin_0			(wallace_cout[6][0] ),
	.cin_1			(wallace_cout[6][1] ),
	.cin_2			(wallace_cout[6][2] ),
	.cin_3			(wallace_cout[6][3] ),
	.cin_4			(wallace_cout[6][4] ),
	.cin_5			(wallace_cout[6][5] ),
	.cin_6			(wallace_cout[6][6] ),
	.cin_7			(wallace_cout[6][7] ),
	.cin_8			(wallace_cout[6][8] ),
	.cin_9			(wallace_cout[6][9] ),
	.cin_10			(wallace_cout[6][10]),
	.cin_11			(wallace_cout[6][11]),
	.cin_12			(wallace_cout[6][12]),
	.cin_13			(wallace_cout[6][13]),
	.cin_14			(wallace_cout[6][14]),
	.cout_0			(wallace_cout[7][0] ),
	.cout_1			(wallace_cout[7][1] ),
	.cout_2			(wallace_cout[7][2] ),
	.cout_3			(wallace_cout[7][3] ),
	.cout_4			(wallace_cout[7][4] ),
	.cout_5			(wallace_cout[7][5] ),
	.cout_6			(wallace_cout[7][6] ),
	.cout_7			(wallace_cout[7][7] ),
	.cout_8			(wallace_cout[7][8] ),
	.cout_9			(wallace_cout[7][9] ),
	.cout_10		(wallace_cout[7][10]),
	.cout_11		(wallace_cout[7][11]),
	.cout_12		(wallace_cout[7][12]),
	.cout_13		(wallace_cout[7][13]),
	.cout_14		(wallace_cout[7][14]),
	.wallace_c		(wallace_c[7]		),
	.wallace_s		(wallace_s[7]		)
);
wallace_tree wallace_tree_8(
	.wallace_input	(wallace_input[8]	),
	.cin_0			(wallace_cout[7][0] ),
	.cin_1			(wallace_cout[7][1] ),
	.cin_2			(wallace_cout[7][2] ),
	.cin_3			(wallace_cout[7][3] ),
	.cin_4			(wallace_cout[7][4] ),
	.cin_5			(wallace_cout[7][5] ),
	.cin_6			(wallace_cout[7][6] ),
	.cin_7			(wallace_cout[7][7] ),
	.cin_8			(wallace_cout[7][8] ),
	.cin_9			(wallace_cout[7][9] ),
	.cin_10			(wallace_cout[7][10]),
	.cin_11			(wallace_cout[7][11]),
	.cin_12			(wallace_cout[7][12]),
	.cin_13			(wallace_cout[7][13]),
	.cin_14			(wallace_cout[7][14]),
	.cout_0			(wallace_cout[8][0] ),
	.cout_1			(wallace_cout[8][1] ),
	.cout_2			(wallace_cout[8][2] ),
	.cout_3			(wallace_cout[8][3] ),
	.cout_4			(wallace_cout[8][4] ),
	.cout_5			(wallace_cout[8][5] ),
	.cout_6			(wallace_cout[8][6] ),
	.cout_7			(wallace_cout[8][7] ),
	.cout_8			(wallace_cout[8][8] ),
	.cout_9			(wallace_cout[8][9] ),
	.cout_10		(wallace_cout[8][10]),
	.cout_11		(wallace_cout[8][11]),
	.cout_12		(wallace_cout[8][12]),
	.cout_13		(wallace_cout[8][13]),
	.cout_14		(wallace_cout[8][14]),
	.wallace_c		(wallace_c[8]		),
	.wallace_s		(wallace_s[8]		)
);
wallace_tree wallace_tree_9(
	.wallace_input	(wallace_input[9]	),
	.cin_0			(wallace_cout[8][0] ),
	.cin_1			(wallace_cout[8][1] ),
	.cin_2			(wallace_cout[8][2] ),
	.cin_3			(wallace_cout[8][3] ),
	.cin_4			(wallace_cout[8][4] ),
	.cin_5			(wallace_cout[8][5] ),
	.cin_6			(wallace_cout[8][6] ),
	.cin_7			(wallace_cout[8][7] ),
	.cin_8			(wallace_cout[8][8] ),
	.cin_9			(wallace_cout[8][9] ),
	.cin_10			(wallace_cout[8][10]),
	.cin_11			(wallace_cout[8][11]),
	.cin_12			(wallace_cout[8][12]),
	.cin_13			(wallace_cout[8][13]),
	.cin_14			(wallace_cout[8][14]),
	.cout_0			(wallace_cout[9][0] ),
	.cout_1			(wallace_cout[9][1] ),
	.cout_2			(wallace_cout[9][2] ),
	.cout_3			(wallace_cout[9][3] ),
	.cout_4			(wallace_cout[9][4] ),
	.cout_5			(wallace_cout[9][5] ),
	.cout_6			(wallace_cout[9][6] ),
	.cout_7			(wallace_cout[9][7] ),
	.cout_8			(wallace_cout[9][8] ),
	.cout_9			(wallace_cout[9][9] ),
	.cout_10		(wallace_cout[9][10]),
	.cout_11		(wallace_cout[9][11]),
	.cout_12		(wallace_cout[9][12]),
	.cout_13		(wallace_cout[9][13]),
	.cout_14		(wallace_cout[9][14]),
	.wallace_c		(wallace_c[9]		),
	.wallace_s		(wallace_s[9]		)
);
wallace_tree wallace_tree_10(
	.wallace_input	(wallace_input[10]	),
	.cin_0			(wallace_cout[9][0] ),
	.cin_1			(wallace_cout[9][1] ),
	.cin_2			(wallace_cout[9][2] ),
	.cin_3			(wallace_cout[9][3] ),
	.cin_4			(wallace_cout[9][4] ),
	.cin_5			(wallace_cout[9][5] ),
	.cin_6			(wallace_cout[9][6] ),
	.cin_7			(wallace_cout[9][7] ),
	.cin_8			(wallace_cout[9][8] ),
	.cin_9			(wallace_cout[9][9] ),
	.cin_10			(wallace_cout[9][10]),
	.cin_11			(wallace_cout[9][11]),
	.cin_12			(wallace_cout[9][12]),
	.cin_13			(wallace_cout[9][13]),
	.cin_14			(wallace_cout[9][14]),
	.cout_0			(wallace_cout[10][0] ),
	.cout_1			(wallace_cout[10][1] ),
	.cout_2			(wallace_cout[10][2] ),
	.cout_3			(wallace_cout[10][3] ),
	.cout_4			(wallace_cout[10][4] ),
	.cout_5			(wallace_cout[10][5] ),
	.cout_6			(wallace_cout[10][6] ),
	.cout_7			(wallace_cout[10][7] ),
	.cout_8			(wallace_cout[10][8] ),
	.cout_9			(wallace_cout[10][9] ),
	.cout_10		(wallace_cout[10][10]),
	.cout_11		(wallace_cout[10][11]),
	.cout_12		(wallace_cout[10][12]),
	.cout_13		(wallace_cout[10][13]),
	.cout_14		(wallace_cout[10][14]),
	.wallace_c		(wallace_c[10]		),
	.wallace_s		(wallace_s[10]		)
);
wallace_tree wallace_tree_11(
	.wallace_input	(wallace_input[11]	),
	.cin_0			(wallace_cout[10][0] ),
	.cin_1			(wallace_cout[10][1] ),
	.cin_2			(wallace_cout[10][2] ),
	.cin_3			(wallace_cout[10][3] ),
	.cin_4			(wallace_cout[10][4] ),
	.cin_5			(wallace_cout[10][5] ),
	.cin_6			(wallace_cout[10][6] ),
	.cin_7			(wallace_cout[10][7] ),
	.cin_8			(wallace_cout[10][8] ),
	.cin_9			(wallace_cout[10][9] ),
	.cin_10			(wallace_cout[10][10]),
	.cin_11			(wallace_cout[10][11]),
	.cin_12			(wallace_cout[10][12]),
	.cin_13			(wallace_cout[10][13]),
	.cin_14			(wallace_cout[10][14]),
	.cout_0			(wallace_cout[11][0] ),
	.cout_1			(wallace_cout[11][1] ),
	.cout_2			(wallace_cout[11][2] ),
	.cout_3			(wallace_cout[11][3] ),
	.cout_4			(wallace_cout[11][4] ),
	.cout_5			(wallace_cout[11][5] ),
	.cout_6			(wallace_cout[11][6] ),
	.cout_7			(wallace_cout[11][7] ),
	.cout_8			(wallace_cout[11][8] ),
	.cout_9			(wallace_cout[11][9] ),
	.cout_10		(wallace_cout[11][10]),
	.cout_11		(wallace_cout[11][11]),
	.cout_12		(wallace_cout[11][12]),
	.cout_13		(wallace_cout[11][13]),
	.cout_14		(wallace_cout[11][14]),
	.wallace_c		(wallace_c[11]		),
	.wallace_s		(wallace_s[11]		)
);
wallace_tree wallace_tree_12(
	.wallace_input	(wallace_input[12]	),
	.cin_0			(wallace_cout[11][0] ),
	.cin_1			(wallace_cout[11][1] ),
	.cin_2			(wallace_cout[11][2] ),
	.cin_3			(wallace_cout[11][3] ),
	.cin_4			(wallace_cout[11][4] ),
	.cin_5			(wallace_cout[11][5] ),
	.cin_6			(wallace_cout[11][6] ),
	.cin_7			(wallace_cout[11][7] ),
	.cin_8			(wallace_cout[11][8] ),
	.cin_9			(wallace_cout[11][9] ),
	.cin_10			(wallace_cout[11][10]),
	.cin_11			(wallace_cout[11][11]),
	.cin_12			(wallace_cout[11][12]),
	.cin_13			(wallace_cout[11][13]),
	.cin_14			(wallace_cout[11][14]),
	.cout_0			(wallace_cout[12][0] ),
	.cout_1			(wallace_cout[12][1] ),
	.cout_2			(wallace_cout[12][2] ),
	.cout_3			(wallace_cout[12][3] ),
	.cout_4			(wallace_cout[12][4] ),
	.cout_5			(wallace_cout[12][5] ),
	.cout_6			(wallace_cout[12][6] ),
	.cout_7			(wallace_cout[12][7] ),
	.cout_8			(wallace_cout[12][8] ),
	.cout_9			(wallace_cout[12][9] ),
	.cout_10		(wallace_cout[12][10]),
	.cout_11		(wallace_cout[12][11]),
	.cout_12		(wallace_cout[12][12]),
	.cout_13		(wallace_cout[12][13]),
	.cout_14		(wallace_cout[12][14]),
	.wallace_c		(wallace_c[12]		),
	.wallace_s		(wallace_s[12]		)
);
wallace_tree wallace_tree_13(
	.wallace_input	(wallace_input[13]	),
	.cin_0			(wallace_cout[12][0] ),
	.cin_1			(wallace_cout[12][1] ),
	.cin_2			(wallace_cout[12][2] ),
	.cin_3			(wallace_cout[12][3] ),
	.cin_4			(wallace_cout[12][4] ),
	.cin_5			(wallace_cout[12][5] ),
	.cin_6			(wallace_cout[12][6] ),
	.cin_7			(wallace_cout[12][7] ),
	.cin_8			(wallace_cout[12][8] ),
	.cin_9			(wallace_cout[12][9] ),
	.cin_10			(wallace_cout[12][10]),
	.cin_11			(wallace_cout[12][11]),
	.cin_12			(wallace_cout[12][12]),
	.cin_13			(wallace_cout[12][13]),
	.cin_14			(wallace_cout[12][14]),
	.cout_0			(wallace_cout[13][0] ),
	.cout_1			(wallace_cout[13][1] ),
	.cout_2			(wallace_cout[13][2] ),
	.cout_3			(wallace_cout[13][3] ),
	.cout_4			(wallace_cout[13][4] ),
	.cout_5			(wallace_cout[13][5] ),
	.cout_6			(wallace_cout[13][6] ),
	.cout_7			(wallace_cout[13][7] ),
	.cout_8			(wallace_cout[13][8] ),
	.cout_9			(wallace_cout[13][9] ),
	.cout_10		(wallace_cout[13][10]),
	.cout_11		(wallace_cout[13][11]),
	.cout_12		(wallace_cout[13][12]),
	.cout_13		(wallace_cout[13][13]),
	.cout_14		(wallace_cout[13][14]),
	.wallace_c		(wallace_c[13]		),
	.wallace_s		(wallace_s[13]		)
);
wallace_tree wallace_tree_14(
	.wallace_input	(wallace_input[14]	),
	.cin_0			(wallace_cout[13][0] ),
	.cin_1			(wallace_cout[13][1] ),
	.cin_2			(wallace_cout[13][2] ),
	.cin_3			(wallace_cout[13][3] ),
	.cin_4			(wallace_cout[13][4] ),
	.cin_5			(wallace_cout[13][5] ),
	.cin_6			(wallace_cout[13][6] ),
	.cin_7			(wallace_cout[13][7] ),
	.cin_8			(wallace_cout[13][8] ),
	.cin_9			(wallace_cout[13][9] ),
	.cin_10			(wallace_cout[13][10]),
	.cin_11			(wallace_cout[13][11]),
	.cin_12			(wallace_cout[13][12]),
	.cin_13			(wallace_cout[13][13]),
	.cin_14			(wallace_cout[13][14]),
	.cout_0			(wallace_cout[14][0] ),
	.cout_1			(wallace_cout[14][1] ),
	.cout_2			(wallace_cout[14][2] ),
	.cout_3			(wallace_cout[14][3] ),
	.cout_4			(wallace_cout[14][4] ),
	.cout_5			(wallace_cout[14][5] ),
	.cout_6			(wallace_cout[14][6] ),
	.cout_7			(wallace_cout[14][7] ),
	.cout_8			(wallace_cout[14][8] ),
	.cout_9			(wallace_cout[14][9] ),
	.cout_10		(wallace_cout[14][10]),
	.cout_11		(wallace_cout[14][11]),
	.cout_12		(wallace_cout[14][12]),
	.cout_13		(wallace_cout[14][13]),
	.cout_14		(wallace_cout[14][14]),
	.wallace_c		(wallace_c[14]		),
	.wallace_s		(wallace_s[14]		)
);
wallace_tree wallace_tree_15(
	.wallace_input	(wallace_input[15]	),
	.cin_0			(wallace_cout[14][0] ),
	.cin_1			(wallace_cout[14][1] ),
	.cin_2			(wallace_cout[14][2] ),
	.cin_3			(wallace_cout[14][3] ),
	.cin_4			(wallace_cout[14][4] ),
	.cin_5			(wallace_cout[14][5] ),
	.cin_6			(wallace_cout[14][6] ),
	.cin_7			(wallace_cout[14][7] ),
	.cin_8			(wallace_cout[14][8] ),
	.cin_9			(wallace_cout[14][9] ),
	.cin_10			(wallace_cout[14][10]),
	.cin_11			(wallace_cout[14][11]),
	.cin_12			(wallace_cout[14][12]),
	.cin_13			(wallace_cout[14][13]),
	.cin_14			(wallace_cout[14][14]),
	.cout_0			(wallace_cout[15][0] ),
	.cout_1			(wallace_cout[15][1] ),
	.cout_2			(wallace_cout[15][2] ),
	.cout_3			(wallace_cout[15][3] ),
	.cout_4			(wallace_cout[15][4] ),
	.cout_5			(wallace_cout[15][5] ),
	.cout_6			(wallace_cout[15][6] ),
	.cout_7			(wallace_cout[15][7] ),
	.cout_8			(wallace_cout[15][8] ),
	.cout_9			(wallace_cout[15][9] ),
	.cout_10		(wallace_cout[15][10]),
	.cout_11		(wallace_cout[15][11]),
	.cout_12		(wallace_cout[15][12]),
	.cout_13		(wallace_cout[15][13]),
	.cout_14		(wallace_cout[15][14]),
	.wallace_c		(wallace_c[15]		),
	.wallace_s		(wallace_s[15]		)
);
wallace_tree wallace_tree_16(
	.wallace_input	(wallace_input[16]	),
	.cin_0			(wallace_cout[15][0] ),
	.cin_1			(wallace_cout[15][1] ),
	.cin_2			(wallace_cout[15][2] ),
	.cin_3			(wallace_cout[15][3] ),
	.cin_4			(wallace_cout[15][4] ),
	.cin_5			(wallace_cout[15][5] ),
	.cin_6			(wallace_cout[15][6] ),
	.cin_7			(wallace_cout[15][7] ),
	.cin_8			(wallace_cout[15][8] ),
	.cin_9			(wallace_cout[15][9] ),
	.cin_10			(wallace_cout[15][10]),
	.cin_11			(wallace_cout[15][11]),
	.cin_12			(wallace_cout[15][12]),
	.cin_13			(wallace_cout[15][13]),
	.cin_14			(wallace_cout[15][14]),
	.cout_0			(wallace_cout[16][0] ),
	.cout_1			(wallace_cout[16][1] ),
	.cout_2			(wallace_cout[16][2] ),
	.cout_3			(wallace_cout[16][3] ),
	.cout_4			(wallace_cout[16][4] ),
	.cout_5			(wallace_cout[16][5] ),
	.cout_6			(wallace_cout[16][6] ),
	.cout_7			(wallace_cout[16][7] ),
	.cout_8			(wallace_cout[16][8] ),
	.cout_9			(wallace_cout[16][9] ),
	.cout_10		(wallace_cout[16][10]),
	.cout_11		(wallace_cout[16][11]),
	.cout_12		(wallace_cout[16][12]),
	.cout_13		(wallace_cout[16][13]),
	.cout_14		(wallace_cout[16][14]),
	.wallace_c		(wallace_c[16]		),
	.wallace_s		(wallace_s[16]		)
);
wallace_tree wallace_tree_17(
	.wallace_input	(wallace_input[17]	),
	.cin_0			(wallace_cout[16][0] ),
	.cin_1			(wallace_cout[16][1] ),
	.cin_2			(wallace_cout[16][2] ),
	.cin_3			(wallace_cout[16][3] ),
	.cin_4			(wallace_cout[16][4] ),
	.cin_5			(wallace_cout[16][5] ),
	.cin_6			(wallace_cout[16][6] ),
	.cin_7			(wallace_cout[16][7] ),
	.cin_8			(wallace_cout[16][8] ),
	.cin_9			(wallace_cout[16][9] ),
	.cin_10			(wallace_cout[16][10]),
	.cin_11			(wallace_cout[16][11]),
	.cin_12			(wallace_cout[16][12]),
	.cin_13			(wallace_cout[16][13]),
	.cin_14			(wallace_cout[16][14]),
	.cout_0			(wallace_cout[17][0] ),
	.cout_1			(wallace_cout[17][1] ),
	.cout_2			(wallace_cout[17][2] ),
	.cout_3			(wallace_cout[17][3] ),
	.cout_4			(wallace_cout[17][4] ),
	.cout_5			(wallace_cout[17][5] ),
	.cout_6			(wallace_cout[17][6] ),
	.cout_7			(wallace_cout[17][7] ),
	.cout_8			(wallace_cout[17][8] ),
	.cout_9			(wallace_cout[17][9] ),
	.cout_10		(wallace_cout[17][10]),
	.cout_11		(wallace_cout[17][11]),
	.cout_12		(wallace_cout[17][12]),
	.cout_13		(wallace_cout[17][13]),
	.cout_14		(wallace_cout[17][14]),
	.wallace_c		(wallace_c[17]		),
	.wallace_s		(wallace_s[17]		)
);
wallace_tree wallace_tree_18(
	.wallace_input	(wallace_input[18]	),
	.cin_0			(wallace_cout[17][0] ),
	.cin_1			(wallace_cout[17][1] ),
	.cin_2			(wallace_cout[17][2] ),
	.cin_3			(wallace_cout[17][3] ),
	.cin_4			(wallace_cout[17][4] ),
	.cin_5			(wallace_cout[17][5] ),
	.cin_6			(wallace_cout[17][6] ),
	.cin_7			(wallace_cout[17][7] ),
	.cin_8			(wallace_cout[17][8] ),
	.cin_9			(wallace_cout[17][9] ),
	.cin_10			(wallace_cout[17][10]),
	.cin_11			(wallace_cout[17][11]),
	.cin_12			(wallace_cout[17][12]),
	.cin_13			(wallace_cout[17][13]),
	.cin_14			(wallace_cout[17][14]),
	.cout_0			(wallace_cout[18][0] ),
	.cout_1			(wallace_cout[18][1] ),
	.cout_2			(wallace_cout[18][2] ),
	.cout_3			(wallace_cout[18][3] ),
	.cout_4			(wallace_cout[18][4] ),
	.cout_5			(wallace_cout[18][5] ),
	.cout_6			(wallace_cout[18][6] ),
	.cout_7			(wallace_cout[18][7] ),
	.cout_8			(wallace_cout[18][8] ),
	.cout_9			(wallace_cout[18][9] ),
	.cout_10		(wallace_cout[18][10]),
	.cout_11		(wallace_cout[18][11]),
	.cout_12		(wallace_cout[18][12]),
	.cout_13		(wallace_cout[18][13]),
	.cout_14		(wallace_cout[18][14]),
	.wallace_c		(wallace_c[18]		),
	.wallace_s		(wallace_s[18]		)
);
wallace_tree wallace_tree_19(
	.wallace_input	(wallace_input[19]	),
	.cin_0			(wallace_cout[18][0] ),
	.cin_1			(wallace_cout[18][1] ),
	.cin_2			(wallace_cout[18][2] ),
	.cin_3			(wallace_cout[18][3] ),
	.cin_4			(wallace_cout[18][4] ),
	.cin_5			(wallace_cout[18][5] ),
	.cin_6			(wallace_cout[18][6] ),
	.cin_7			(wallace_cout[18][7] ),
	.cin_8			(wallace_cout[18][8] ),
	.cin_9			(wallace_cout[18][9] ),
	.cin_10			(wallace_cout[18][10]),
	.cin_11			(wallace_cout[18][11]),
	.cin_12			(wallace_cout[18][12]),
	.cin_13			(wallace_cout[18][13]),
	.cin_14			(wallace_cout[18][14]),
	.cout_0			(wallace_cout[19][0] ),
	.cout_1			(wallace_cout[19][1] ),
	.cout_2			(wallace_cout[19][2] ),
	.cout_3			(wallace_cout[19][3] ),
	.cout_4			(wallace_cout[19][4] ),
	.cout_5			(wallace_cout[19][5] ),
	.cout_6			(wallace_cout[19][6] ),
	.cout_7			(wallace_cout[19][7] ),
	.cout_8			(wallace_cout[19][8] ),
	.cout_9			(wallace_cout[19][9] ),
	.cout_10		(wallace_cout[19][10]),
	.cout_11		(wallace_cout[19][11]),
	.cout_12		(wallace_cout[19][12]),
	.cout_13		(wallace_cout[19][13]),
	.cout_14		(wallace_cout[19][14]),
	.wallace_c		(wallace_c[19]		),
	.wallace_s		(wallace_s[19]		)
);
wallace_tree wallace_tree_20(
	.wallace_input	(wallace_input[20]	),
	.cin_0			(wallace_cout[19][0] ),
	.cin_1			(wallace_cout[19][1] ),
	.cin_2			(wallace_cout[19][2] ),
	.cin_3			(wallace_cout[19][3] ),
	.cin_4			(wallace_cout[19][4] ),
	.cin_5			(wallace_cout[19][5] ),
	.cin_6			(wallace_cout[19][6] ),
	.cin_7			(wallace_cout[19][7] ),
	.cin_8			(wallace_cout[19][8] ),
	.cin_9			(wallace_cout[19][9] ),
	.cin_10			(wallace_cout[19][10]),
	.cin_11			(wallace_cout[19][11]),
	.cin_12			(wallace_cout[19][12]),
	.cin_13			(wallace_cout[19][13]),
	.cin_14			(wallace_cout[19][14]),
	.cout_0			(wallace_cout[20][0] ),
	.cout_1			(wallace_cout[20][1] ),
	.cout_2			(wallace_cout[20][2] ),
	.cout_3			(wallace_cout[20][3] ),
	.cout_4			(wallace_cout[20][4] ),
	.cout_5			(wallace_cout[20][5] ),
	.cout_6			(wallace_cout[20][6] ),
	.cout_7			(wallace_cout[20][7] ),
	.cout_8			(wallace_cout[20][8] ),
	.cout_9			(wallace_cout[20][9] ),
	.cout_10		(wallace_cout[20][10]),
	.cout_11		(wallace_cout[20][11]),
	.cout_12		(wallace_cout[20][12]),
	.cout_13		(wallace_cout[20][13]),
	.cout_14		(wallace_cout[20][14]),
	.wallace_c		(wallace_c[20]		),
	.wallace_s		(wallace_s[20]		)
);
wallace_tree wallace_tree_21(
	.wallace_input	(wallace_input[21]	),
	.cin_0			(wallace_cout[20][0] ),
	.cin_1			(wallace_cout[20][1] ),
	.cin_2			(wallace_cout[20][2] ),
	.cin_3			(wallace_cout[20][3] ),
	.cin_4			(wallace_cout[20][4] ),
	.cin_5			(wallace_cout[20][5] ),
	.cin_6			(wallace_cout[20][6] ),
	.cin_7			(wallace_cout[20][7] ),
	.cin_8			(wallace_cout[20][8] ),
	.cin_9			(wallace_cout[20][9] ),
	.cin_10			(wallace_cout[20][10]),
	.cin_11			(wallace_cout[20][11]),
	.cin_12			(wallace_cout[20][12]),
	.cin_13			(wallace_cout[20][13]),
	.cin_14			(wallace_cout[20][14]),
	.cout_0			(wallace_cout[21][0] ),
	.cout_1			(wallace_cout[21][1] ),
	.cout_2			(wallace_cout[21][2] ),
	.cout_3			(wallace_cout[21][3] ),
	.cout_4			(wallace_cout[21][4] ),
	.cout_5			(wallace_cout[21][5] ),
	.cout_6			(wallace_cout[21][6] ),
	.cout_7			(wallace_cout[21][7] ),
	.cout_8			(wallace_cout[21][8] ),
	.cout_9			(wallace_cout[21][9] ),
	.cout_10		(wallace_cout[21][10]),
	.cout_11		(wallace_cout[21][11]),
	.cout_12		(wallace_cout[21][12]),
	.cout_13		(wallace_cout[21][13]),
	.cout_14		(wallace_cout[21][14]),
	.wallace_c		(wallace_c[21]		),
	.wallace_s		(wallace_s[21]		)
);
wallace_tree wallace_tree_22(
	.wallace_input	(wallace_input[22]	),
	.cin_0			(wallace_cout[21][0] ),
	.cin_1			(wallace_cout[21][1] ),
	.cin_2			(wallace_cout[21][2] ),
	.cin_3			(wallace_cout[21][3] ),
	.cin_4			(wallace_cout[21][4] ),
	.cin_5			(wallace_cout[21][5] ),
	.cin_6			(wallace_cout[21][6] ),
	.cin_7			(wallace_cout[21][7] ),
	.cin_8			(wallace_cout[21][8] ),
	.cin_9			(wallace_cout[21][9] ),
	.cin_10			(wallace_cout[21][10]),
	.cin_11			(wallace_cout[21][11]),
	.cin_12			(wallace_cout[21][12]),
	.cin_13			(wallace_cout[21][13]),
	.cin_14			(wallace_cout[21][14]),
	.cout_0			(wallace_cout[22][0] ),
	.cout_1			(wallace_cout[22][1] ),
	.cout_2			(wallace_cout[22][2] ),
	.cout_3			(wallace_cout[22][3] ),
	.cout_4			(wallace_cout[22][4] ),
	.cout_5			(wallace_cout[22][5] ),
	.cout_6			(wallace_cout[22][6] ),
	.cout_7			(wallace_cout[22][7] ),
	.cout_8			(wallace_cout[22][8] ),
	.cout_9			(wallace_cout[22][9] ),
	.cout_10		(wallace_cout[22][10]),
	.cout_11		(wallace_cout[22][11]),
	.cout_12		(wallace_cout[22][12]),
	.cout_13		(wallace_cout[22][13]),
	.cout_14		(wallace_cout[22][14]),
	.wallace_c		(wallace_c[22]		),
	.wallace_s		(wallace_s[22]		)
);
wallace_tree wallace_tree_23(
	.wallace_input	(wallace_input[23]	),
	.cin_0			(wallace_cout[22][0] ),
	.cin_1			(wallace_cout[22][1] ),
	.cin_2			(wallace_cout[22][2] ),
	.cin_3			(wallace_cout[22][3] ),
	.cin_4			(wallace_cout[22][4] ),
	.cin_5			(wallace_cout[22][5] ),
	.cin_6			(wallace_cout[22][6] ),
	.cin_7			(wallace_cout[22][7] ),
	.cin_8			(wallace_cout[22][8] ),
	.cin_9			(wallace_cout[22][9] ),
	.cin_10			(wallace_cout[22][10]),
	.cin_11			(wallace_cout[22][11]),
	.cin_12			(wallace_cout[22][12]),
	.cin_13			(wallace_cout[22][13]),
	.cin_14			(wallace_cout[22][14]),
	.cout_0			(wallace_cout[23][0] ),
	.cout_1			(wallace_cout[23][1] ),
	.cout_2			(wallace_cout[23][2] ),
	.cout_3			(wallace_cout[23][3] ),
	.cout_4			(wallace_cout[23][4] ),
	.cout_5			(wallace_cout[23][5] ),
	.cout_6			(wallace_cout[23][6] ),
	.cout_7			(wallace_cout[23][7] ),
	.cout_8			(wallace_cout[23][8] ),
	.cout_9			(wallace_cout[23][9] ),
	.cout_10		(wallace_cout[23][10]),
	.cout_11		(wallace_cout[23][11]),
	.cout_12		(wallace_cout[23][12]),
	.cout_13		(wallace_cout[23][13]),
	.cout_14		(wallace_cout[23][14]),
	.wallace_c		(wallace_c[23]		),
	.wallace_s		(wallace_s[23]		)
);
wallace_tree wallace_tree_24(
	.wallace_input	(wallace_input[24]	),
	.cin_0			(wallace_cout[23][0] ),
	.cin_1			(wallace_cout[23][1] ),
	.cin_2			(wallace_cout[23][2] ),
	.cin_3			(wallace_cout[23][3] ),
	.cin_4			(wallace_cout[23][4] ),
	.cin_5			(wallace_cout[23][5] ),
	.cin_6			(wallace_cout[23][6] ),
	.cin_7			(wallace_cout[23][7] ),
	.cin_8			(wallace_cout[23][8] ),
	.cin_9			(wallace_cout[23][9] ),
	.cin_10			(wallace_cout[23][10]),
	.cin_11			(wallace_cout[23][11]),
	.cin_12			(wallace_cout[23][12]),
	.cin_13			(wallace_cout[23][13]),
	.cin_14			(wallace_cout[23][14]),
	.cout_0			(wallace_cout[24][0] ),
	.cout_1			(wallace_cout[24][1] ),
	.cout_2			(wallace_cout[24][2] ),
	.cout_3			(wallace_cout[24][3] ),
	.cout_4			(wallace_cout[24][4] ),
	.cout_5			(wallace_cout[24][5] ),
	.cout_6			(wallace_cout[24][6] ),
	.cout_7			(wallace_cout[24][7] ),
	.cout_8			(wallace_cout[24][8] ),
	.cout_9			(wallace_cout[24][9] ),
	.cout_10		(wallace_cout[24][10]),
	.cout_11		(wallace_cout[24][11]),
	.cout_12		(wallace_cout[24][12]),
	.cout_13		(wallace_cout[24][13]),
	.cout_14		(wallace_cout[24][14]),
	.wallace_c		(wallace_c[24]		),
	.wallace_s		(wallace_s[24]		)
);
wallace_tree wallace_tree_25(
	.wallace_input	(wallace_input[25]	),
	.cin_0			(wallace_cout[24][0] ),
	.cin_1			(wallace_cout[24][1] ),
	.cin_2			(wallace_cout[24][2] ),
	.cin_3			(wallace_cout[24][3] ),
	.cin_4			(wallace_cout[24][4] ),
	.cin_5			(wallace_cout[24][5] ),
	.cin_6			(wallace_cout[24][6] ),
	.cin_7			(wallace_cout[24][7] ),
	.cin_8			(wallace_cout[24][8] ),
	.cin_9			(wallace_cout[24][9] ),
	.cin_10			(wallace_cout[24][10]),
	.cin_11			(wallace_cout[24][11]),
	.cin_12			(wallace_cout[24][12]),
	.cin_13			(wallace_cout[24][13]),
	.cin_14			(wallace_cout[24][14]),
	.cout_0			(wallace_cout[25][0] ),
	.cout_1			(wallace_cout[25][1] ),
	.cout_2			(wallace_cout[25][2] ),
	.cout_3			(wallace_cout[25][3] ),
	.cout_4			(wallace_cout[25][4] ),
	.cout_5			(wallace_cout[25][5] ),
	.cout_6			(wallace_cout[25][6] ),
	.cout_7			(wallace_cout[25][7] ),
	.cout_8			(wallace_cout[25][8] ),
	.cout_9			(wallace_cout[25][9] ),
	.cout_10		(wallace_cout[25][10]),
	.cout_11		(wallace_cout[25][11]),
	.cout_12		(wallace_cout[25][12]),
	.cout_13		(wallace_cout[25][13]),
	.cout_14		(wallace_cout[25][14]),
	.wallace_c		(wallace_c[25]		),
	.wallace_s		(wallace_s[25]		)
);
wallace_tree wallace_tree_26(
	.wallace_input	(wallace_input[26]	),
	.cin_0			(wallace_cout[25][0] ),
	.cin_1			(wallace_cout[25][1] ),
	.cin_2			(wallace_cout[25][2] ),
	.cin_3			(wallace_cout[25][3] ),
	.cin_4			(wallace_cout[25][4] ),
	.cin_5			(wallace_cout[25][5] ),
	.cin_6			(wallace_cout[25][6] ),
	.cin_7			(wallace_cout[25][7] ),
	.cin_8			(wallace_cout[25][8] ),
	.cin_9			(wallace_cout[25][9] ),
	.cin_10			(wallace_cout[25][10]),
	.cin_11			(wallace_cout[25][11]),
	.cin_12			(wallace_cout[25][12]),
	.cin_13			(wallace_cout[25][13]),
	.cin_14			(wallace_cout[25][14]),
	.cout_0			(wallace_cout[26][0] ),
	.cout_1			(wallace_cout[26][1] ),
	.cout_2			(wallace_cout[26][2] ),
	.cout_3			(wallace_cout[26][3] ),
	.cout_4			(wallace_cout[26][4] ),
	.cout_5			(wallace_cout[26][5] ),
	.cout_6			(wallace_cout[26][6] ),
	.cout_7			(wallace_cout[26][7] ),
	.cout_8			(wallace_cout[26][8] ),
	.cout_9			(wallace_cout[26][9] ),
	.cout_10		(wallace_cout[26][10]),
	.cout_11		(wallace_cout[26][11]),
	.cout_12		(wallace_cout[26][12]),
	.cout_13		(wallace_cout[26][13]),
	.cout_14		(wallace_cout[26][14]),
	.wallace_c		(wallace_c[26]		),
	.wallace_s		(wallace_s[26]		)
);
wallace_tree wallace_tree_27(
	.wallace_input	(wallace_input[27]	),
	.cin_0			(wallace_cout[26][0] ),
	.cin_1			(wallace_cout[26][1] ),
	.cin_2			(wallace_cout[26][2] ),
	.cin_3			(wallace_cout[26][3] ),
	.cin_4			(wallace_cout[26][4] ),
	.cin_5			(wallace_cout[26][5] ),
	.cin_6			(wallace_cout[26][6] ),
	.cin_7			(wallace_cout[26][7] ),
	.cin_8			(wallace_cout[26][8] ),
	.cin_9			(wallace_cout[26][9] ),
	.cin_10			(wallace_cout[26][10]),
	.cin_11			(wallace_cout[26][11]),
	.cin_12			(wallace_cout[26][12]),
	.cin_13			(wallace_cout[26][13]),
	.cin_14			(wallace_cout[26][14]),
	.cout_0			(wallace_cout[27][0] ),
	.cout_1			(wallace_cout[27][1] ),
	.cout_2			(wallace_cout[27][2] ),
	.cout_3			(wallace_cout[27][3] ),
	.cout_4			(wallace_cout[27][4] ),
	.cout_5			(wallace_cout[27][5] ),
	.cout_6			(wallace_cout[27][6] ),
	.cout_7			(wallace_cout[27][7] ),
	.cout_8			(wallace_cout[27][8] ),
	.cout_9			(wallace_cout[27][9] ),
	.cout_10		(wallace_cout[27][10]),
	.cout_11		(wallace_cout[27][11]),
	.cout_12		(wallace_cout[27][12]),
	.cout_13		(wallace_cout[27][13]),
	.cout_14		(wallace_cout[27][14]),
	.wallace_c		(wallace_c[27]		),
	.wallace_s		(wallace_s[27]		)
);
wallace_tree wallace_tree_28(
	.wallace_input	(wallace_input[28]	),
	.cin_0			(wallace_cout[27][0] ),
	.cin_1			(wallace_cout[27][1] ),
	.cin_2			(wallace_cout[27][2] ),
	.cin_3			(wallace_cout[27][3] ),
	.cin_4			(wallace_cout[27][4] ),
	.cin_5			(wallace_cout[27][5] ),
	.cin_6			(wallace_cout[27][6] ),
	.cin_7			(wallace_cout[27][7] ),
	.cin_8			(wallace_cout[27][8] ),
	.cin_9			(wallace_cout[27][9] ),
	.cin_10			(wallace_cout[27][10]),
	.cin_11			(wallace_cout[27][11]),
	.cin_12			(wallace_cout[27][12]),
	.cin_13			(wallace_cout[27][13]),
	.cin_14			(wallace_cout[27][14]),
	.cout_0			(wallace_cout[28][0] ),
	.cout_1			(wallace_cout[28][1] ),
	.cout_2			(wallace_cout[28][2] ),
	.cout_3			(wallace_cout[28][3] ),
	.cout_4			(wallace_cout[28][4] ),
	.cout_5			(wallace_cout[28][5] ),
	.cout_6			(wallace_cout[28][6] ),
	.cout_7			(wallace_cout[28][7] ),
	.cout_8			(wallace_cout[28][8] ),
	.cout_9			(wallace_cout[28][9] ),
	.cout_10		(wallace_cout[28][10]),
	.cout_11		(wallace_cout[28][11]),
	.cout_12		(wallace_cout[28][12]),
	.cout_13		(wallace_cout[28][13]),
	.cout_14		(wallace_cout[28][14]),
	.wallace_c		(wallace_c[28]		),
	.wallace_s		(wallace_s[28]		)
);
wallace_tree wallace_tree_29(
	.wallace_input	(wallace_input[29]	),
	.cin_0			(wallace_cout[28][0] ),
	.cin_1			(wallace_cout[28][1] ),
	.cin_2			(wallace_cout[28][2] ),
	.cin_3			(wallace_cout[28][3] ),
	.cin_4			(wallace_cout[28][4] ),
	.cin_5			(wallace_cout[28][5] ),
	.cin_6			(wallace_cout[28][6] ),
	.cin_7			(wallace_cout[28][7] ),
	.cin_8			(wallace_cout[28][8] ),
	.cin_9			(wallace_cout[28][9] ),
	.cin_10			(wallace_cout[28][10]),
	.cin_11			(wallace_cout[28][11]),
	.cin_12			(wallace_cout[28][12]),
	.cin_13			(wallace_cout[28][13]),
	.cin_14			(wallace_cout[28][14]),
	.cout_0			(wallace_cout[29][0] ),
	.cout_1			(wallace_cout[29][1] ),
	.cout_2			(wallace_cout[29][2] ),
	.cout_3			(wallace_cout[29][3] ),
	.cout_4			(wallace_cout[29][4] ),
	.cout_5			(wallace_cout[29][5] ),
	.cout_6			(wallace_cout[29][6] ),
	.cout_7			(wallace_cout[29][7] ),
	.cout_8			(wallace_cout[29][8] ),
	.cout_9			(wallace_cout[29][9] ),
	.cout_10		(wallace_cout[29][10]),
	.cout_11		(wallace_cout[29][11]),
	.cout_12		(wallace_cout[29][12]),
	.cout_13		(wallace_cout[29][13]),
	.cout_14		(wallace_cout[29][14]),
	.wallace_c		(wallace_c[29]		),
	.wallace_s		(wallace_s[29]		)
);
wallace_tree wallace_tree_30(
	.wallace_input	(wallace_input[30]	),
	.cin_0			(wallace_cout[29][0] ),
	.cin_1			(wallace_cout[29][1] ),
	.cin_2			(wallace_cout[29][2] ),
	.cin_3			(wallace_cout[29][3] ),
	.cin_4			(wallace_cout[29][4] ),
	.cin_5			(wallace_cout[29][5] ),
	.cin_6			(wallace_cout[29][6] ),
	.cin_7			(wallace_cout[29][7] ),
	.cin_8			(wallace_cout[29][8] ),
	.cin_9			(wallace_cout[29][9] ),
	.cin_10			(wallace_cout[29][10]),
	.cin_11			(wallace_cout[29][11]),
	.cin_12			(wallace_cout[29][12]),
	.cin_13			(wallace_cout[29][13]),
	.cin_14			(wallace_cout[29][14]),
	.cout_0			(wallace_cout[30][0] ),
	.cout_1			(wallace_cout[30][1] ),
	.cout_2			(wallace_cout[30][2] ),
	.cout_3			(wallace_cout[30][3] ),
	.cout_4			(wallace_cout[30][4] ),
	.cout_5			(wallace_cout[30][5] ),
	.cout_6			(wallace_cout[30][6] ),
	.cout_7			(wallace_cout[30][7] ),
	.cout_8			(wallace_cout[30][8] ),
	.cout_9			(wallace_cout[30][9] ),
	.cout_10		(wallace_cout[30][10]),
	.cout_11		(wallace_cout[30][11]),
	.cout_12		(wallace_cout[30][12]),
	.cout_13		(wallace_cout[30][13]),
	.cout_14		(wallace_cout[30][14]),
	.wallace_c		(wallace_c[30]		),
	.wallace_s		(wallace_s[30]		)
);
wallace_tree wallace_tree_31(
	.wallace_input	(wallace_input[31]	),
	.cin_0			(wallace_cout[30][0] ),
	.cin_1			(wallace_cout[30][1] ),
	.cin_2			(wallace_cout[30][2] ),
	.cin_3			(wallace_cout[30][3] ),
	.cin_4			(wallace_cout[30][4] ),
	.cin_5			(wallace_cout[30][5] ),
	.cin_6			(wallace_cout[30][6] ),
	.cin_7			(wallace_cout[30][7] ),
	.cin_8			(wallace_cout[30][8] ),
	.cin_9			(wallace_cout[30][9] ),
	.cin_10			(wallace_cout[30][10]),
	.cin_11			(wallace_cout[30][11]),
	.cin_12			(wallace_cout[30][12]),
	.cin_13			(wallace_cout[30][13]),
	.cin_14			(wallace_cout[30][14]),
	.cout_0			(wallace_cout[31][0] ),
	.cout_1			(wallace_cout[31][1] ),
	.cout_2			(wallace_cout[31][2] ),
	.cout_3			(wallace_cout[31][3] ),
	.cout_4			(wallace_cout[31][4] ),
	.cout_5			(wallace_cout[31][5] ),
	.cout_6			(wallace_cout[31][6] ),
	.cout_7			(wallace_cout[31][7] ),
	.cout_8			(wallace_cout[31][8] ),
	.cout_9			(wallace_cout[31][9] ),
	.cout_10		(wallace_cout[31][10]),
	.cout_11		(wallace_cout[31][11]),
	.cout_12		(wallace_cout[31][12]),
	.cout_13		(wallace_cout[31][13]),
	.cout_14		(wallace_cout[31][14]),
	.wallace_c		(wallace_c[31]		),
	.wallace_s		(wallace_s[31]		)
);
wallace_tree wallace_tree_32(
	.wallace_input	(wallace_input[32]	),
	.cin_0			(wallace_cout[31][0] ),
	.cin_1			(wallace_cout[31][1] ),
	.cin_2			(wallace_cout[31][2] ),
	.cin_3			(wallace_cout[31][3] ),
	.cin_4			(wallace_cout[31][4] ),
	.cin_5			(wallace_cout[31][5] ),
	.cin_6			(wallace_cout[31][6] ),
	.cin_7			(wallace_cout[31][7] ),
	.cin_8			(wallace_cout[31][8] ),
	.cin_9			(wallace_cout[31][9] ),
	.cin_10			(wallace_cout[31][10]),
	.cin_11			(wallace_cout[31][11]),
	.cin_12			(wallace_cout[31][12]),
	.cin_13			(wallace_cout[31][13]),
	.cin_14			(wallace_cout[31][14]),
	.cout_0			(wallace_cout[32][0] ),
	.cout_1			(wallace_cout[32][1] ),
	.cout_2			(wallace_cout[32][2] ),
	.cout_3			(wallace_cout[32][3] ),
	.cout_4			(wallace_cout[32][4] ),
	.cout_5			(wallace_cout[32][5] ),
	.cout_6			(wallace_cout[32][6] ),
	.cout_7			(wallace_cout[32][7] ),
	.cout_8			(wallace_cout[32][8] ),
	.cout_9			(wallace_cout[32][9] ),
	.cout_10		(wallace_cout[32][10]),
	.cout_11		(wallace_cout[32][11]),
	.cout_12		(wallace_cout[32][12]),
	.cout_13		(wallace_cout[32][13]),
	.cout_14		(wallace_cout[32][14]),
	.wallace_c		(wallace_c[32]		),
	.wallace_s		(wallace_s[32]		)
);
wallace_tree wallace_tree_33(
	.wallace_input	(wallace_input[33]	),
	.cin_0			(wallace_cout[32][0] ),
	.cin_1			(wallace_cout[32][1] ),
	.cin_2			(wallace_cout[32][2] ),
	.cin_3			(wallace_cout[32][3] ),
	.cin_4			(wallace_cout[32][4] ),
	.cin_5			(wallace_cout[32][5] ),
	.cin_6			(wallace_cout[32][6] ),
	.cin_7			(wallace_cout[32][7] ),
	.cin_8			(wallace_cout[32][8] ),
	.cin_9			(wallace_cout[32][9] ),
	.cin_10			(wallace_cout[32][10]),
	.cin_11			(wallace_cout[32][11]),
	.cin_12			(wallace_cout[32][12]),
	.cin_13			(wallace_cout[32][13]),
	.cin_14			(wallace_cout[32][14]),
	.cout_0			(wallace_cout[33][0] ),
	.cout_1			(wallace_cout[33][1] ),
	.cout_2			(wallace_cout[33][2] ),
	.cout_3			(wallace_cout[33][3] ),
	.cout_4			(wallace_cout[33][4] ),
	.cout_5			(wallace_cout[33][5] ),
	.cout_6			(wallace_cout[33][6] ),
	.cout_7			(wallace_cout[33][7] ),
	.cout_8			(wallace_cout[33][8] ),
	.cout_9			(wallace_cout[33][9] ),
	.cout_10		(wallace_cout[33][10]),
	.cout_11		(wallace_cout[33][11]),
	.cout_12		(wallace_cout[33][12]),
	.cout_13		(wallace_cout[33][13]),
	.cout_14		(wallace_cout[33][14]),
	.wallace_c		(wallace_c[33]		),
	.wallace_s		(wallace_s[33]		)
);
wallace_tree wallace_tree_34(
	.wallace_input	(wallace_input[34]	),
	.cin_0			(wallace_cout[33][0] ),
	.cin_1			(wallace_cout[33][1] ),
	.cin_2			(wallace_cout[33][2] ),
	.cin_3			(wallace_cout[33][3] ),
	.cin_4			(wallace_cout[33][4] ),
	.cin_5			(wallace_cout[33][5] ),
	.cin_6			(wallace_cout[33][6] ),
	.cin_7			(wallace_cout[33][7] ),
	.cin_8			(wallace_cout[33][8] ),
	.cin_9			(wallace_cout[33][9] ),
	.cin_10			(wallace_cout[33][10]),
	.cin_11			(wallace_cout[33][11]),
	.cin_12			(wallace_cout[33][12]),
	.cin_13			(wallace_cout[33][13]),
	.cin_14			(wallace_cout[33][14]),
	.cout_0			(wallace_cout[34][0] ),
	.cout_1			(wallace_cout[34][1] ),
	.cout_2			(wallace_cout[34][2] ),
	.cout_3			(wallace_cout[34][3] ),
	.cout_4			(wallace_cout[34][4] ),
	.cout_5			(wallace_cout[34][5] ),
	.cout_6			(wallace_cout[34][6] ),
	.cout_7			(wallace_cout[34][7] ),
	.cout_8			(wallace_cout[34][8] ),
	.cout_9			(wallace_cout[34][9] ),
	.cout_10		(wallace_cout[34][10]),
	.cout_11		(wallace_cout[34][11]),
	.cout_12		(wallace_cout[34][12]),
	.cout_13		(wallace_cout[34][13]),
	.cout_14		(wallace_cout[34][14]),
	.wallace_c		(wallace_c[34]		),
	.wallace_s		(wallace_s[34]		)
);
wallace_tree wallace_tree_35(
	.wallace_input	(wallace_input[35]	),
	.cin_0			(wallace_cout[34][0] ),
	.cin_1			(wallace_cout[34][1] ),
	.cin_2			(wallace_cout[34][2] ),
	.cin_3			(wallace_cout[34][3] ),
	.cin_4			(wallace_cout[34][4] ),
	.cin_5			(wallace_cout[34][5] ),
	.cin_6			(wallace_cout[34][6] ),
	.cin_7			(wallace_cout[34][7] ),
	.cin_8			(wallace_cout[34][8] ),
	.cin_9			(wallace_cout[34][9] ),
	.cin_10			(wallace_cout[34][10]),
	.cin_11			(wallace_cout[34][11]),
	.cin_12			(wallace_cout[34][12]),
	.cin_13			(wallace_cout[34][13]),
	.cin_14			(wallace_cout[34][14]),
	.cout_0			(wallace_cout[35][0] ),
	.cout_1			(wallace_cout[35][1] ),
	.cout_2			(wallace_cout[35][2] ),
	.cout_3			(wallace_cout[35][3] ),
	.cout_4			(wallace_cout[35][4] ),
	.cout_5			(wallace_cout[35][5] ),
	.cout_6			(wallace_cout[35][6] ),
	.cout_7			(wallace_cout[35][7] ),
	.cout_8			(wallace_cout[35][8] ),
	.cout_9			(wallace_cout[35][9] ),
	.cout_10		(wallace_cout[35][10]),
	.cout_11		(wallace_cout[35][11]),
	.cout_12		(wallace_cout[35][12]),
	.cout_13		(wallace_cout[35][13]),
	.cout_14		(wallace_cout[35][14]),
	.wallace_c		(wallace_c[35]		),
	.wallace_s		(wallace_s[35]		)
);
wallace_tree wallace_tree_36(
	.wallace_input	(wallace_input[36]	),
	.cin_0			(wallace_cout[35][0] ),
	.cin_1			(wallace_cout[35][1] ),
	.cin_2			(wallace_cout[35][2] ),
	.cin_3			(wallace_cout[35][3] ),
	.cin_4			(wallace_cout[35][4] ),
	.cin_5			(wallace_cout[35][5] ),
	.cin_6			(wallace_cout[35][6] ),
	.cin_7			(wallace_cout[35][7] ),
	.cin_8			(wallace_cout[35][8] ),
	.cin_9			(wallace_cout[35][9] ),
	.cin_10			(wallace_cout[35][10]),
	.cin_11			(wallace_cout[35][11]),
	.cin_12			(wallace_cout[35][12]),
	.cin_13			(wallace_cout[35][13]),
	.cin_14			(wallace_cout[35][14]),
	.cout_0			(wallace_cout[36][0] ),
	.cout_1			(wallace_cout[36][1] ),
	.cout_2			(wallace_cout[36][2] ),
	.cout_3			(wallace_cout[36][3] ),
	.cout_4			(wallace_cout[36][4] ),
	.cout_5			(wallace_cout[36][5] ),
	.cout_6			(wallace_cout[36][6] ),
	.cout_7			(wallace_cout[36][7] ),
	.cout_8			(wallace_cout[36][8] ),
	.cout_9			(wallace_cout[36][9] ),
	.cout_10		(wallace_cout[36][10]),
	.cout_11		(wallace_cout[36][11]),
	.cout_12		(wallace_cout[36][12]),
	.cout_13		(wallace_cout[36][13]),
	.cout_14		(wallace_cout[36][14]),
	.wallace_c		(wallace_c[36]		),
	.wallace_s		(wallace_s[36]		)
);
wallace_tree wallace_tree_37(
	.wallace_input	(wallace_input[37]	),
	.cin_0			(wallace_cout[36][0] ),
	.cin_1			(wallace_cout[36][1] ),
	.cin_2			(wallace_cout[36][2] ),
	.cin_3			(wallace_cout[36][3] ),
	.cin_4			(wallace_cout[36][4] ),
	.cin_5			(wallace_cout[36][5] ),
	.cin_6			(wallace_cout[36][6] ),
	.cin_7			(wallace_cout[36][7] ),
	.cin_8			(wallace_cout[36][8] ),
	.cin_9			(wallace_cout[36][9] ),
	.cin_10			(wallace_cout[36][10]),
	.cin_11			(wallace_cout[36][11]),
	.cin_12			(wallace_cout[36][12]),
	.cin_13			(wallace_cout[36][13]),
	.cin_14			(wallace_cout[36][14]),
	.cout_0			(wallace_cout[37][0] ),
	.cout_1			(wallace_cout[37][1] ),
	.cout_2			(wallace_cout[37][2] ),
	.cout_3			(wallace_cout[37][3] ),
	.cout_4			(wallace_cout[37][4] ),
	.cout_5			(wallace_cout[37][5] ),
	.cout_6			(wallace_cout[37][6] ),
	.cout_7			(wallace_cout[37][7] ),
	.cout_8			(wallace_cout[37][8] ),
	.cout_9			(wallace_cout[37][9] ),
	.cout_10		(wallace_cout[37][10]),
	.cout_11		(wallace_cout[37][11]),
	.cout_12		(wallace_cout[37][12]),
	.cout_13		(wallace_cout[37][13]),
	.cout_14		(wallace_cout[37][14]),
	.wallace_c		(wallace_c[37]		),
	.wallace_s		(wallace_s[37]		)
);
wallace_tree wallace_tree_38(
	.wallace_input	(wallace_input[38]	),
	.cin_0			(wallace_cout[37][0] ),
	.cin_1			(wallace_cout[37][1] ),
	.cin_2			(wallace_cout[37][2] ),
	.cin_3			(wallace_cout[37][3] ),
	.cin_4			(wallace_cout[37][4] ),
	.cin_5			(wallace_cout[37][5] ),
	.cin_6			(wallace_cout[37][6] ),
	.cin_7			(wallace_cout[37][7] ),
	.cin_8			(wallace_cout[37][8] ),
	.cin_9			(wallace_cout[37][9] ),
	.cin_10			(wallace_cout[37][10]),
	.cin_11			(wallace_cout[37][11]),
	.cin_12			(wallace_cout[37][12]),
	.cin_13			(wallace_cout[37][13]),
	.cin_14			(wallace_cout[37][14]),
	.cout_0			(wallace_cout[38][0] ),
	.cout_1			(wallace_cout[38][1] ),
	.cout_2			(wallace_cout[38][2] ),
	.cout_3			(wallace_cout[38][3] ),
	.cout_4			(wallace_cout[38][4] ),
	.cout_5			(wallace_cout[38][5] ),
	.cout_6			(wallace_cout[38][6] ),
	.cout_7			(wallace_cout[38][7] ),
	.cout_8			(wallace_cout[38][8] ),
	.cout_9			(wallace_cout[38][9] ),
	.cout_10		(wallace_cout[38][10]),
	.cout_11		(wallace_cout[38][11]),
	.cout_12		(wallace_cout[38][12]),
	.cout_13		(wallace_cout[38][13]),
	.cout_14		(wallace_cout[38][14]),
	.wallace_c		(wallace_c[38]		),
	.wallace_s		(wallace_s[38]		)
);
wallace_tree wallace_tree_39(
	.wallace_input	(wallace_input[39]	),
	.cin_0			(wallace_cout[38][0] ),
	.cin_1			(wallace_cout[38][1] ),
	.cin_2			(wallace_cout[38][2] ),
	.cin_3			(wallace_cout[38][3] ),
	.cin_4			(wallace_cout[38][4] ),
	.cin_5			(wallace_cout[38][5] ),
	.cin_6			(wallace_cout[38][6] ),
	.cin_7			(wallace_cout[38][7] ),
	.cin_8			(wallace_cout[38][8] ),
	.cin_9			(wallace_cout[38][9] ),
	.cin_10			(wallace_cout[38][10]),
	.cin_11			(wallace_cout[38][11]),
	.cin_12			(wallace_cout[38][12]),
	.cin_13			(wallace_cout[38][13]),
	.cin_14			(wallace_cout[38][14]),
	.cout_0			(wallace_cout[39][0] ),
	.cout_1			(wallace_cout[39][1] ),
	.cout_2			(wallace_cout[39][2] ),
	.cout_3			(wallace_cout[39][3] ),
	.cout_4			(wallace_cout[39][4] ),
	.cout_5			(wallace_cout[39][5] ),
	.cout_6			(wallace_cout[39][6] ),
	.cout_7			(wallace_cout[39][7] ),
	.cout_8			(wallace_cout[39][8] ),
	.cout_9			(wallace_cout[39][9] ),
	.cout_10		(wallace_cout[39][10]),
	.cout_11		(wallace_cout[39][11]),
	.cout_12		(wallace_cout[39][12]),
	.cout_13		(wallace_cout[39][13]),
	.cout_14		(wallace_cout[39][14]),
	.wallace_c		(wallace_c[39]		),
	.wallace_s		(wallace_s[39]		)
);
wallace_tree wallace_tree_40(
	.wallace_input	(wallace_input[40]	),
	.cin_0			(wallace_cout[39][0] ),
	.cin_1			(wallace_cout[39][1] ),
	.cin_2			(wallace_cout[39][2] ),
	.cin_3			(wallace_cout[39][3] ),
	.cin_4			(wallace_cout[39][4] ),
	.cin_5			(wallace_cout[39][5] ),
	.cin_6			(wallace_cout[39][6] ),
	.cin_7			(wallace_cout[39][7] ),
	.cin_8			(wallace_cout[39][8] ),
	.cin_9			(wallace_cout[39][9] ),
	.cin_10			(wallace_cout[39][10]),
	.cin_11			(wallace_cout[39][11]),
	.cin_12			(wallace_cout[39][12]),
	.cin_13			(wallace_cout[39][13]),
	.cin_14			(wallace_cout[39][14]),
	.cout_0			(wallace_cout[40][0] ),
	.cout_1			(wallace_cout[40][1] ),
	.cout_2			(wallace_cout[40][2] ),
	.cout_3			(wallace_cout[40][3] ),
	.cout_4			(wallace_cout[40][4] ),
	.cout_5			(wallace_cout[40][5] ),
	.cout_6			(wallace_cout[40][6] ),
	.cout_7			(wallace_cout[40][7] ),
	.cout_8			(wallace_cout[40][8] ),
	.cout_9			(wallace_cout[40][9] ),
	.cout_10		(wallace_cout[40][10]),
	.cout_11		(wallace_cout[40][11]),
	.cout_12		(wallace_cout[40][12]),
	.cout_13		(wallace_cout[40][13]),
	.cout_14		(wallace_cout[40][14]),
	.wallace_c		(wallace_c[40]		),
	.wallace_s		(wallace_s[40]		)
);
wallace_tree wallace_tree_41(
	.wallace_input	(wallace_input[41]	),
	.cin_0			(wallace_cout[40][0] ),
	.cin_1			(wallace_cout[40][1] ),
	.cin_2			(wallace_cout[40][2] ),
	.cin_3			(wallace_cout[40][3] ),
	.cin_4			(wallace_cout[40][4] ),
	.cin_5			(wallace_cout[40][5] ),
	.cin_6			(wallace_cout[40][6] ),
	.cin_7			(wallace_cout[40][7] ),
	.cin_8			(wallace_cout[40][8] ),
	.cin_9			(wallace_cout[40][9] ),
	.cin_10			(wallace_cout[40][10]),
	.cin_11			(wallace_cout[40][11]),
	.cin_12			(wallace_cout[40][12]),
	.cin_13			(wallace_cout[40][13]),
	.cin_14			(wallace_cout[40][14]),
	.cout_0			(wallace_cout[41][0] ),
	.cout_1			(wallace_cout[41][1] ),
	.cout_2			(wallace_cout[41][2] ),
	.cout_3			(wallace_cout[41][3] ),
	.cout_4			(wallace_cout[41][4] ),
	.cout_5			(wallace_cout[41][5] ),
	.cout_6			(wallace_cout[41][6] ),
	.cout_7			(wallace_cout[41][7] ),
	.cout_8			(wallace_cout[41][8] ),
	.cout_9			(wallace_cout[41][9] ),
	.cout_10		(wallace_cout[41][10]),
	.cout_11		(wallace_cout[41][11]),
	.cout_12		(wallace_cout[41][12]),
	.cout_13		(wallace_cout[41][13]),
	.cout_14		(wallace_cout[41][14]),
	.wallace_c		(wallace_c[41]		),
	.wallace_s		(wallace_s[41]		)
);
wallace_tree wallace_tree_42(
	.wallace_input	(wallace_input[42]	),
	.cin_0			(wallace_cout[41][0] ),
	.cin_1			(wallace_cout[41][1] ),
	.cin_2			(wallace_cout[41][2] ),
	.cin_3			(wallace_cout[41][3] ),
	.cin_4			(wallace_cout[41][4] ),
	.cin_5			(wallace_cout[41][5] ),
	.cin_6			(wallace_cout[41][6] ),
	.cin_7			(wallace_cout[41][7] ),
	.cin_8			(wallace_cout[41][8] ),
	.cin_9			(wallace_cout[41][9] ),
	.cin_10			(wallace_cout[41][10]),
	.cin_11			(wallace_cout[41][11]),
	.cin_12			(wallace_cout[41][12]),
	.cin_13			(wallace_cout[41][13]),
	.cin_14			(wallace_cout[41][14]),
	.cout_0			(wallace_cout[42][0] ),
	.cout_1			(wallace_cout[42][1] ),
	.cout_2			(wallace_cout[42][2] ),
	.cout_3			(wallace_cout[42][3] ),
	.cout_4			(wallace_cout[42][4] ),
	.cout_5			(wallace_cout[42][5] ),
	.cout_6			(wallace_cout[42][6] ),
	.cout_7			(wallace_cout[42][7] ),
	.cout_8			(wallace_cout[42][8] ),
	.cout_9			(wallace_cout[42][9] ),
	.cout_10		(wallace_cout[42][10]),
	.cout_11		(wallace_cout[42][11]),
	.cout_12		(wallace_cout[42][12]),
	.cout_13		(wallace_cout[42][13]),
	.cout_14		(wallace_cout[42][14]),
	.wallace_c		(wallace_c[42]		),
	.wallace_s		(wallace_s[42]		)
);
wallace_tree wallace_tree_43(
	.wallace_input	(wallace_input[43]	),
	.cin_0			(wallace_cout[42][0] ),
	.cin_1			(wallace_cout[42][1] ),
	.cin_2			(wallace_cout[42][2] ),
	.cin_3			(wallace_cout[42][3] ),
	.cin_4			(wallace_cout[42][4] ),
	.cin_5			(wallace_cout[42][5] ),
	.cin_6			(wallace_cout[42][6] ),
	.cin_7			(wallace_cout[42][7] ),
	.cin_8			(wallace_cout[42][8] ),
	.cin_9			(wallace_cout[42][9] ),
	.cin_10			(wallace_cout[42][10]),
	.cin_11			(wallace_cout[42][11]),
	.cin_12			(wallace_cout[42][12]),
	.cin_13			(wallace_cout[42][13]),
	.cin_14			(wallace_cout[42][14]),
	.cout_0			(wallace_cout[43][0] ),
	.cout_1			(wallace_cout[43][1] ),
	.cout_2			(wallace_cout[43][2] ),
	.cout_3			(wallace_cout[43][3] ),
	.cout_4			(wallace_cout[43][4] ),
	.cout_5			(wallace_cout[43][5] ),
	.cout_6			(wallace_cout[43][6] ),
	.cout_7			(wallace_cout[43][7] ),
	.cout_8			(wallace_cout[43][8] ),
	.cout_9			(wallace_cout[43][9] ),
	.cout_10		(wallace_cout[43][10]),
	.cout_11		(wallace_cout[43][11]),
	.cout_12		(wallace_cout[43][12]),
	.cout_13		(wallace_cout[43][13]),
	.cout_14		(wallace_cout[43][14]),
	.wallace_c		(wallace_c[43]		),
	.wallace_s		(wallace_s[43]		)
);
wallace_tree wallace_tree_44(
	.wallace_input	(wallace_input[44]	),
	.cin_0			(wallace_cout[43][0] ),
	.cin_1			(wallace_cout[43][1] ),
	.cin_2			(wallace_cout[43][2] ),
	.cin_3			(wallace_cout[43][3] ),
	.cin_4			(wallace_cout[43][4] ),
	.cin_5			(wallace_cout[43][5] ),
	.cin_6			(wallace_cout[43][6] ),
	.cin_7			(wallace_cout[43][7] ),
	.cin_8			(wallace_cout[43][8] ),
	.cin_9			(wallace_cout[43][9] ),
	.cin_10			(wallace_cout[43][10]),
	.cin_11			(wallace_cout[43][11]),
	.cin_12			(wallace_cout[43][12]),
	.cin_13			(wallace_cout[43][13]),
	.cin_14			(wallace_cout[43][14]),
	.cout_0			(wallace_cout[44][0] ),
	.cout_1			(wallace_cout[44][1] ),
	.cout_2			(wallace_cout[44][2] ),
	.cout_3			(wallace_cout[44][3] ),
	.cout_4			(wallace_cout[44][4] ),
	.cout_5			(wallace_cout[44][5] ),
	.cout_6			(wallace_cout[44][6] ),
	.cout_7			(wallace_cout[44][7] ),
	.cout_8			(wallace_cout[44][8] ),
	.cout_9			(wallace_cout[44][9] ),
	.cout_10		(wallace_cout[44][10]),
	.cout_11		(wallace_cout[44][11]),
	.cout_12		(wallace_cout[44][12]),
	.cout_13		(wallace_cout[44][13]),
	.cout_14		(wallace_cout[44][14]),
	.wallace_c		(wallace_c[44]		),
	.wallace_s		(wallace_s[44]		)
);
wallace_tree wallace_tree_45(
	.wallace_input	(wallace_input[45]	),
	.cin_0			(wallace_cout[44][0] ),
	.cin_1			(wallace_cout[44][1] ),
	.cin_2			(wallace_cout[44][2] ),
	.cin_3			(wallace_cout[44][3] ),
	.cin_4			(wallace_cout[44][4] ),
	.cin_5			(wallace_cout[44][5] ),
	.cin_6			(wallace_cout[44][6] ),
	.cin_7			(wallace_cout[44][7] ),
	.cin_8			(wallace_cout[44][8] ),
	.cin_9			(wallace_cout[44][9] ),
	.cin_10			(wallace_cout[44][10]),
	.cin_11			(wallace_cout[44][11]),
	.cin_12			(wallace_cout[44][12]),
	.cin_13			(wallace_cout[44][13]),
	.cin_14			(wallace_cout[44][14]),
	.cout_0			(wallace_cout[45][0] ),
	.cout_1			(wallace_cout[45][1] ),
	.cout_2			(wallace_cout[45][2] ),
	.cout_3			(wallace_cout[45][3] ),
	.cout_4			(wallace_cout[45][4] ),
	.cout_5			(wallace_cout[45][5] ),
	.cout_6			(wallace_cout[45][6] ),
	.cout_7			(wallace_cout[45][7] ),
	.cout_8			(wallace_cout[45][8] ),
	.cout_9			(wallace_cout[45][9] ),
	.cout_10		(wallace_cout[45][10]),
	.cout_11		(wallace_cout[45][11]),
	.cout_12		(wallace_cout[45][12]),
	.cout_13		(wallace_cout[45][13]),
	.cout_14		(wallace_cout[45][14]),
	.wallace_c		(wallace_c[45]		),
	.wallace_s		(wallace_s[45]		)
);
wallace_tree wallace_tree_46(
	.wallace_input	(wallace_input[46]	),
	.cin_0			(wallace_cout[45][0] ),
	.cin_1			(wallace_cout[45][1] ),
	.cin_2			(wallace_cout[45][2] ),
	.cin_3			(wallace_cout[45][3] ),
	.cin_4			(wallace_cout[45][4] ),
	.cin_5			(wallace_cout[45][5] ),
	.cin_6			(wallace_cout[45][6] ),
	.cin_7			(wallace_cout[45][7] ),
	.cin_8			(wallace_cout[45][8] ),
	.cin_9			(wallace_cout[45][9] ),
	.cin_10			(wallace_cout[45][10]),
	.cin_11			(wallace_cout[45][11]),
	.cin_12			(wallace_cout[45][12]),
	.cin_13			(wallace_cout[45][13]),
	.cin_14			(wallace_cout[45][14]),
	.cout_0			(wallace_cout[46][0] ),
	.cout_1			(wallace_cout[46][1] ),
	.cout_2			(wallace_cout[46][2] ),
	.cout_3			(wallace_cout[46][3] ),
	.cout_4			(wallace_cout[46][4] ),
	.cout_5			(wallace_cout[46][5] ),
	.cout_6			(wallace_cout[46][6] ),
	.cout_7			(wallace_cout[46][7] ),
	.cout_8			(wallace_cout[46][8] ),
	.cout_9			(wallace_cout[46][9] ),
	.cout_10		(wallace_cout[46][10]),
	.cout_11		(wallace_cout[46][11]),
	.cout_12		(wallace_cout[46][12]),
	.cout_13		(wallace_cout[46][13]),
	.cout_14		(wallace_cout[46][14]),
	.wallace_c		(wallace_c[46]		),
	.wallace_s		(wallace_s[46]		)
);
wallace_tree wallace_tree_47(
	.wallace_input	(wallace_input[47]	),
	.cin_0			(wallace_cout[46][0] ),
	.cin_1			(wallace_cout[46][1] ),
	.cin_2			(wallace_cout[46][2] ),
	.cin_3			(wallace_cout[46][3] ),
	.cin_4			(wallace_cout[46][4] ),
	.cin_5			(wallace_cout[46][5] ),
	.cin_6			(wallace_cout[46][6] ),
	.cin_7			(wallace_cout[46][7] ),
	.cin_8			(wallace_cout[46][8] ),
	.cin_9			(wallace_cout[46][9] ),
	.cin_10			(wallace_cout[46][10]),
	.cin_11			(wallace_cout[46][11]),
	.cin_12			(wallace_cout[46][12]),
	.cin_13			(wallace_cout[46][13]),
	.cin_14			(wallace_cout[46][14]),
	.cout_0			(wallace_cout[47][0] ),
	.cout_1			(wallace_cout[47][1] ),
	.cout_2			(wallace_cout[47][2] ),
	.cout_3			(wallace_cout[47][3] ),
	.cout_4			(wallace_cout[47][4] ),
	.cout_5			(wallace_cout[47][5] ),
	.cout_6			(wallace_cout[47][6] ),
	.cout_7			(wallace_cout[47][7] ),
	.cout_8			(wallace_cout[47][8] ),
	.cout_9			(wallace_cout[47][9] ),
	.cout_10		(wallace_cout[47][10]),
	.cout_11		(wallace_cout[47][11]),
	.cout_12		(wallace_cout[47][12]),
	.cout_13		(wallace_cout[47][13]),
	.cout_14		(wallace_cout[47][14]),
	.wallace_c		(wallace_c[47]		),
	.wallace_s		(wallace_s[47]		)
);
wallace_tree wallace_tree_48(
	.wallace_input	(wallace_input[48]	),
	.cin_0			(wallace_cout[47][0] ),
	.cin_1			(wallace_cout[47][1] ),
	.cin_2			(wallace_cout[47][2] ),
	.cin_3			(wallace_cout[47][3] ),
	.cin_4			(wallace_cout[47][4] ),
	.cin_5			(wallace_cout[47][5] ),
	.cin_6			(wallace_cout[47][6] ),
	.cin_7			(wallace_cout[47][7] ),
	.cin_8			(wallace_cout[47][8] ),
	.cin_9			(wallace_cout[47][9] ),
	.cin_10			(wallace_cout[47][10]),
	.cin_11			(wallace_cout[47][11]),
	.cin_12			(wallace_cout[47][12]),
	.cin_13			(wallace_cout[47][13]),
	.cin_14			(wallace_cout[47][14]),
	.cout_0			(wallace_cout[48][0] ),
	.cout_1			(wallace_cout[48][1] ),
	.cout_2			(wallace_cout[48][2] ),
	.cout_3			(wallace_cout[48][3] ),
	.cout_4			(wallace_cout[48][4] ),
	.cout_5			(wallace_cout[48][5] ),
	.cout_6			(wallace_cout[48][6] ),
	.cout_7			(wallace_cout[48][7] ),
	.cout_8			(wallace_cout[48][8] ),
	.cout_9			(wallace_cout[48][9] ),
	.cout_10		(wallace_cout[48][10]),
	.cout_11		(wallace_cout[48][11]),
	.cout_12		(wallace_cout[48][12]),
	.cout_13		(wallace_cout[48][13]),
	.cout_14		(wallace_cout[48][14]),
	.wallace_c		(wallace_c[48]		),
	.wallace_s		(wallace_s[48]		)
);
wallace_tree wallace_tree_49(
	.wallace_input	(wallace_input[49]	),
	.cin_0			(wallace_cout[48][0] ),
	.cin_1			(wallace_cout[48][1] ),
	.cin_2			(wallace_cout[48][2] ),
	.cin_3			(wallace_cout[48][3] ),
	.cin_4			(wallace_cout[48][4] ),
	.cin_5			(wallace_cout[48][5] ),
	.cin_6			(wallace_cout[48][6] ),
	.cin_7			(wallace_cout[48][7] ),
	.cin_8			(wallace_cout[48][8] ),
	.cin_9			(wallace_cout[48][9] ),
	.cin_10			(wallace_cout[48][10]),
	.cin_11			(wallace_cout[48][11]),
	.cin_12			(wallace_cout[48][12]),
	.cin_13			(wallace_cout[48][13]),
	.cin_14			(wallace_cout[48][14]),
	.cout_0			(wallace_cout[49][0] ),
	.cout_1			(wallace_cout[49][1] ),
	.cout_2			(wallace_cout[49][2] ),
	.cout_3			(wallace_cout[49][3] ),
	.cout_4			(wallace_cout[49][4] ),
	.cout_5			(wallace_cout[49][5] ),
	.cout_6			(wallace_cout[49][6] ),
	.cout_7			(wallace_cout[49][7] ),
	.cout_8			(wallace_cout[49][8] ),
	.cout_9			(wallace_cout[49][9] ),
	.cout_10		(wallace_cout[49][10]),
	.cout_11		(wallace_cout[49][11]),
	.cout_12		(wallace_cout[49][12]),
	.cout_13		(wallace_cout[49][13]),
	.cout_14		(wallace_cout[49][14]),
	.wallace_c		(wallace_c[49]		),
	.wallace_s		(wallace_s[49]		)
);
wallace_tree wallace_tree_50(
	.wallace_input	(wallace_input[50]	),
	.cin_0			(wallace_cout[49][0] ),
	.cin_1			(wallace_cout[49][1] ),
	.cin_2			(wallace_cout[49][2] ),
	.cin_3			(wallace_cout[49][3] ),
	.cin_4			(wallace_cout[49][4] ),
	.cin_5			(wallace_cout[49][5] ),
	.cin_6			(wallace_cout[49][6] ),
	.cin_7			(wallace_cout[49][7] ),
	.cin_8			(wallace_cout[49][8] ),
	.cin_9			(wallace_cout[49][9] ),
	.cin_10			(wallace_cout[49][10]),
	.cin_11			(wallace_cout[49][11]),
	.cin_12			(wallace_cout[49][12]),
	.cin_13			(wallace_cout[49][13]),
	.cin_14			(wallace_cout[49][14]),
	.cout_0			(wallace_cout[50][0] ),
	.cout_1			(wallace_cout[50][1] ),
	.cout_2			(wallace_cout[50][2] ),
	.cout_3			(wallace_cout[50][3] ),
	.cout_4			(wallace_cout[50][4] ),
	.cout_5			(wallace_cout[50][5] ),
	.cout_6			(wallace_cout[50][6] ),
	.cout_7			(wallace_cout[50][7] ),
	.cout_8			(wallace_cout[50][8] ),
	.cout_9			(wallace_cout[50][9] ),
	.cout_10		(wallace_cout[50][10]),
	.cout_11		(wallace_cout[50][11]),
	.cout_12		(wallace_cout[50][12]),
	.cout_13		(wallace_cout[50][13]),
	.cout_14		(wallace_cout[50][14]),
	.wallace_c		(wallace_c[50]		),
	.wallace_s		(wallace_s[50]		)
);
wallace_tree wallace_tree_51(
	.wallace_input	(wallace_input[51]	),
	.cin_0			(wallace_cout[50][0] ),
	.cin_1			(wallace_cout[50][1] ),
	.cin_2			(wallace_cout[50][2] ),
	.cin_3			(wallace_cout[50][3] ),
	.cin_4			(wallace_cout[50][4] ),
	.cin_5			(wallace_cout[50][5] ),
	.cin_6			(wallace_cout[50][6] ),
	.cin_7			(wallace_cout[50][7] ),
	.cin_8			(wallace_cout[50][8] ),
	.cin_9			(wallace_cout[50][9] ),
	.cin_10			(wallace_cout[50][10]),
	.cin_11			(wallace_cout[50][11]),
	.cin_12			(wallace_cout[50][12]),
	.cin_13			(wallace_cout[50][13]),
	.cin_14			(wallace_cout[50][14]),
	.cout_0			(wallace_cout[51][0] ),
	.cout_1			(wallace_cout[51][1] ),
	.cout_2			(wallace_cout[51][2] ),
	.cout_3			(wallace_cout[51][3] ),
	.cout_4			(wallace_cout[51][4] ),
	.cout_5			(wallace_cout[51][5] ),
	.cout_6			(wallace_cout[51][6] ),
	.cout_7			(wallace_cout[51][7] ),
	.cout_8			(wallace_cout[51][8] ),
	.cout_9			(wallace_cout[51][9] ),
	.cout_10		(wallace_cout[51][10]),
	.cout_11		(wallace_cout[51][11]),
	.cout_12		(wallace_cout[51][12]),
	.cout_13		(wallace_cout[51][13]),
	.cout_14		(wallace_cout[51][14]),
	.wallace_c		(wallace_c[51]		),
	.wallace_s		(wallace_s[51]		)
);
wallace_tree wallace_tree_52(
	.wallace_input	(wallace_input[52]	),
	.cin_0			(wallace_cout[51][0] ),
	.cin_1			(wallace_cout[51][1] ),
	.cin_2			(wallace_cout[51][2] ),
	.cin_3			(wallace_cout[51][3] ),
	.cin_4			(wallace_cout[51][4] ),
	.cin_5			(wallace_cout[51][5] ),
	.cin_6			(wallace_cout[51][6] ),
	.cin_7			(wallace_cout[51][7] ),
	.cin_8			(wallace_cout[51][8] ),
	.cin_9			(wallace_cout[51][9] ),
	.cin_10			(wallace_cout[51][10]),
	.cin_11			(wallace_cout[51][11]),
	.cin_12			(wallace_cout[51][12]),
	.cin_13			(wallace_cout[51][13]),
	.cin_14			(wallace_cout[51][14]),
	.cout_0			(wallace_cout[52][0] ),
	.cout_1			(wallace_cout[52][1] ),
	.cout_2			(wallace_cout[52][2] ),
	.cout_3			(wallace_cout[52][3] ),
	.cout_4			(wallace_cout[52][4] ),
	.cout_5			(wallace_cout[52][5] ),
	.cout_6			(wallace_cout[52][6] ),
	.cout_7			(wallace_cout[52][7] ),
	.cout_8			(wallace_cout[52][8] ),
	.cout_9			(wallace_cout[52][9] ),
	.cout_10		(wallace_cout[52][10]),
	.cout_11		(wallace_cout[52][11]),
	.cout_12		(wallace_cout[52][12]),
	.cout_13		(wallace_cout[52][13]),
	.cout_14		(wallace_cout[52][14]),
	.wallace_c		(wallace_c[52]		),
	.wallace_s		(wallace_s[52]		)
);
wallace_tree wallace_tree_53(
	.wallace_input	(wallace_input[53]	),
	.cin_0			(wallace_cout[52][0] ),
	.cin_1			(wallace_cout[52][1] ),
	.cin_2			(wallace_cout[52][2] ),
	.cin_3			(wallace_cout[52][3] ),
	.cin_4			(wallace_cout[52][4] ),
	.cin_5			(wallace_cout[52][5] ),
	.cin_6			(wallace_cout[52][6] ),
	.cin_7			(wallace_cout[52][7] ),
	.cin_8			(wallace_cout[52][8] ),
	.cin_9			(wallace_cout[52][9] ),
	.cin_10			(wallace_cout[52][10]),
	.cin_11			(wallace_cout[52][11]),
	.cin_12			(wallace_cout[52][12]),
	.cin_13			(wallace_cout[52][13]),
	.cin_14			(wallace_cout[52][14]),
	.cout_0			(wallace_cout[53][0] ),
	.cout_1			(wallace_cout[53][1] ),
	.cout_2			(wallace_cout[53][2] ),
	.cout_3			(wallace_cout[53][3] ),
	.cout_4			(wallace_cout[53][4] ),
	.cout_5			(wallace_cout[53][5] ),
	.cout_6			(wallace_cout[53][6] ),
	.cout_7			(wallace_cout[53][7] ),
	.cout_8			(wallace_cout[53][8] ),
	.cout_9			(wallace_cout[53][9] ),
	.cout_10		(wallace_cout[53][10]),
	.cout_11		(wallace_cout[53][11]),
	.cout_12		(wallace_cout[53][12]),
	.cout_13		(wallace_cout[53][13]),
	.cout_14		(wallace_cout[53][14]),
	.wallace_c		(wallace_c[53]		),
	.wallace_s		(wallace_s[53]		)
);
wallace_tree wallace_tree_54(
	.wallace_input	(wallace_input[54]	),
	.cin_0			(wallace_cout[53][0] ),
	.cin_1			(wallace_cout[53][1] ),
	.cin_2			(wallace_cout[53][2] ),
	.cin_3			(wallace_cout[53][3] ),
	.cin_4			(wallace_cout[53][4] ),
	.cin_5			(wallace_cout[53][5] ),
	.cin_6			(wallace_cout[53][6] ),
	.cin_7			(wallace_cout[53][7] ),
	.cin_8			(wallace_cout[53][8] ),
	.cin_9			(wallace_cout[53][9] ),
	.cin_10			(wallace_cout[53][10]),
	.cin_11			(wallace_cout[53][11]),
	.cin_12			(wallace_cout[53][12]),
	.cin_13			(wallace_cout[53][13]),
	.cin_14			(wallace_cout[53][14]),
	.cout_0			(wallace_cout[54][0] ),
	.cout_1			(wallace_cout[54][1] ),
	.cout_2			(wallace_cout[54][2] ),
	.cout_3			(wallace_cout[54][3] ),
	.cout_4			(wallace_cout[54][4] ),
	.cout_5			(wallace_cout[54][5] ),
	.cout_6			(wallace_cout[54][6] ),
	.cout_7			(wallace_cout[54][7] ),
	.cout_8			(wallace_cout[54][8] ),
	.cout_9			(wallace_cout[54][9] ),
	.cout_10		(wallace_cout[54][10]),
	.cout_11		(wallace_cout[54][11]),
	.cout_12		(wallace_cout[54][12]),
	.cout_13		(wallace_cout[54][13]),
	.cout_14		(wallace_cout[54][14]),
	.wallace_c		(wallace_c[54]		),
	.wallace_s		(wallace_s[54]		)
);
wallace_tree wallace_tree_55(
	.wallace_input	(wallace_input[55]	),
	.cin_0			(wallace_cout[54][0] ),
	.cin_1			(wallace_cout[54][1] ),
	.cin_2			(wallace_cout[54][2] ),
	.cin_3			(wallace_cout[54][3] ),
	.cin_4			(wallace_cout[54][4] ),
	.cin_5			(wallace_cout[54][5] ),
	.cin_6			(wallace_cout[54][6] ),
	.cin_7			(wallace_cout[54][7] ),
	.cin_8			(wallace_cout[54][8] ),
	.cin_9			(wallace_cout[54][9] ),
	.cin_10			(wallace_cout[54][10]),
	.cin_11			(wallace_cout[54][11]),
	.cin_12			(wallace_cout[54][12]),
	.cin_13			(wallace_cout[54][13]),
	.cin_14			(wallace_cout[54][14]),
	.cout_0			(wallace_cout[55][0] ),
	.cout_1			(wallace_cout[55][1] ),
	.cout_2			(wallace_cout[55][2] ),
	.cout_3			(wallace_cout[55][3] ),
	.cout_4			(wallace_cout[55][4] ),
	.cout_5			(wallace_cout[55][5] ),
	.cout_6			(wallace_cout[55][6] ),
	.cout_7			(wallace_cout[55][7] ),
	.cout_8			(wallace_cout[55][8] ),
	.cout_9			(wallace_cout[55][9] ),
	.cout_10		(wallace_cout[55][10]),
	.cout_11		(wallace_cout[55][11]),
	.cout_12		(wallace_cout[55][12]),
	.cout_13		(wallace_cout[55][13]),
	.cout_14		(wallace_cout[55][14]),
	.wallace_c		(wallace_c[55]		),
	.wallace_s		(wallace_s[55]		)
);
wallace_tree wallace_tree_56(
	.wallace_input	(wallace_input[56]	),
	.cin_0			(wallace_cout[55][0] ),
	.cin_1			(wallace_cout[55][1] ),
	.cin_2			(wallace_cout[55][2] ),
	.cin_3			(wallace_cout[55][3] ),
	.cin_4			(wallace_cout[55][4] ),
	.cin_5			(wallace_cout[55][5] ),
	.cin_6			(wallace_cout[55][6] ),
	.cin_7			(wallace_cout[55][7] ),
	.cin_8			(wallace_cout[55][8] ),
	.cin_9			(wallace_cout[55][9] ),
	.cin_10			(wallace_cout[55][10]),
	.cin_11			(wallace_cout[55][11]),
	.cin_12			(wallace_cout[55][12]),
	.cin_13			(wallace_cout[55][13]),
	.cin_14			(wallace_cout[55][14]),
	.cout_0			(wallace_cout[56][0] ),
	.cout_1			(wallace_cout[56][1] ),
	.cout_2			(wallace_cout[56][2] ),
	.cout_3			(wallace_cout[56][3] ),
	.cout_4			(wallace_cout[56][4] ),
	.cout_5			(wallace_cout[56][5] ),
	.cout_6			(wallace_cout[56][6] ),
	.cout_7			(wallace_cout[56][7] ),
	.cout_8			(wallace_cout[56][8] ),
	.cout_9			(wallace_cout[56][9] ),
	.cout_10		(wallace_cout[56][10]),
	.cout_11		(wallace_cout[56][11]),
	.cout_12		(wallace_cout[56][12]),
	.cout_13		(wallace_cout[56][13]),
	.cout_14		(wallace_cout[56][14]),
	.wallace_c		(wallace_c[56]		),
	.wallace_s		(wallace_s[56]		)
);
wallace_tree wallace_tree_57(
	.wallace_input	(wallace_input[57]	),
	.cin_0			(wallace_cout[56][0] ),
	.cin_1			(wallace_cout[56][1] ),
	.cin_2			(wallace_cout[56][2] ),
	.cin_3			(wallace_cout[56][3] ),
	.cin_4			(wallace_cout[56][4] ),
	.cin_5			(wallace_cout[56][5] ),
	.cin_6			(wallace_cout[56][6] ),
	.cin_7			(wallace_cout[56][7] ),
	.cin_8			(wallace_cout[56][8] ),
	.cin_9			(wallace_cout[56][9] ),
	.cin_10			(wallace_cout[56][10]),
	.cin_11			(wallace_cout[56][11]),
	.cin_12			(wallace_cout[56][12]),
	.cin_13			(wallace_cout[56][13]),
	.cin_14			(wallace_cout[56][14]),
	.cout_0			(wallace_cout[57][0] ),
	.cout_1			(wallace_cout[57][1] ),
	.cout_2			(wallace_cout[57][2] ),
	.cout_3			(wallace_cout[57][3] ),
	.cout_4			(wallace_cout[57][4] ),
	.cout_5			(wallace_cout[57][5] ),
	.cout_6			(wallace_cout[57][6] ),
	.cout_7			(wallace_cout[57][7] ),
	.cout_8			(wallace_cout[57][8] ),
	.cout_9			(wallace_cout[57][9] ),
	.cout_10		(wallace_cout[57][10]),
	.cout_11		(wallace_cout[57][11]),
	.cout_12		(wallace_cout[57][12]),
	.cout_13		(wallace_cout[57][13]),
	.cout_14		(wallace_cout[57][14]),
	.wallace_c		(wallace_c[57]		),
	.wallace_s		(wallace_s[57]		)
);
wallace_tree wallace_tree_58(
	.wallace_input	(wallace_input[58]	),
	.cin_0			(wallace_cout[57][0] ),
	.cin_1			(wallace_cout[57][1] ),
	.cin_2			(wallace_cout[57][2] ),
	.cin_3			(wallace_cout[57][3] ),
	.cin_4			(wallace_cout[57][4] ),
	.cin_5			(wallace_cout[57][5] ),
	.cin_6			(wallace_cout[57][6] ),
	.cin_7			(wallace_cout[57][7] ),
	.cin_8			(wallace_cout[57][8] ),
	.cin_9			(wallace_cout[57][9] ),
	.cin_10			(wallace_cout[57][10]),
	.cin_11			(wallace_cout[57][11]),
	.cin_12			(wallace_cout[57][12]),
	.cin_13			(wallace_cout[57][13]),
	.cin_14			(wallace_cout[57][14]),
	.cout_0			(wallace_cout[58][0] ),
	.cout_1			(wallace_cout[58][1] ),
	.cout_2			(wallace_cout[58][2] ),
	.cout_3			(wallace_cout[58][3] ),
	.cout_4			(wallace_cout[58][4] ),
	.cout_5			(wallace_cout[58][5] ),
	.cout_6			(wallace_cout[58][6] ),
	.cout_7			(wallace_cout[58][7] ),
	.cout_8			(wallace_cout[58][8] ),
	.cout_9			(wallace_cout[58][9] ),
	.cout_10		(wallace_cout[58][10]),
	.cout_11		(wallace_cout[58][11]),
	.cout_12		(wallace_cout[58][12]),
	.cout_13		(wallace_cout[58][13]),
	.cout_14		(wallace_cout[58][14]),
	.wallace_c		(wallace_c[58]		),
	.wallace_s		(wallace_s[58]		)
);
wallace_tree wallace_tree_59(
	.wallace_input	(wallace_input[59]   ),
	.cin_0			(wallace_cout[58][0] ),
	.cin_1			(wallace_cout[58][1] ),
	.cin_2			(wallace_cout[58][2] ),
	.cin_3			(wallace_cout[58][3] ),
	.cin_4			(wallace_cout[58][4] ),
	.cin_5			(wallace_cout[58][5] ),
	.cin_6			(wallace_cout[58][6] ),
	.cin_7			(wallace_cout[58][7] ),
	.cin_8			(wallace_cout[58][8] ),
	.cin_9			(wallace_cout[58][9] ),
	.cin_10			(wallace_cout[58][10]),
	.cin_11			(wallace_cout[58][11]),
	.cin_12			(wallace_cout[58][12]),
	.cin_13			(wallace_cout[58][13]),
	.cin_14			(wallace_cout[58][14]),
	.cout_0			(wallace_cout[59][0] ),
	.cout_1			(wallace_cout[59][1] ),
	.cout_2			(wallace_cout[59][2] ),
	.cout_3			(wallace_cout[59][3] ),
	.cout_4			(wallace_cout[59][4] ),
	.cout_5			(wallace_cout[59][5] ),
	.cout_6			(wallace_cout[59][6] ),
	.cout_7			(wallace_cout[59][7] ),
	.cout_8			(wallace_cout[59][8] ),
	.cout_9			(wallace_cout[59][9] ),
	.cout_10		(wallace_cout[59][10]),
	.cout_11		(wallace_cout[59][11]),
	.cout_12		(wallace_cout[59][12]),
	.cout_13		(wallace_cout[59][13]),
	.cout_14		(wallace_cout[59][14]),
	.wallace_c		(wallace_c[59]       ),
	.wallace_s		(wallace_s[59]       )
);
wallace_tree wallace_tree_60(
	.wallace_input	(wallace_input[60]   ),
	.cin_0			(wallace_cout[59][0] ),
	.cin_1			(wallace_cout[59][1] ),
	.cin_2			(wallace_cout[59][2] ),
	.cin_3			(wallace_cout[59][3] ),
	.cin_4			(wallace_cout[59][4] ),
	.cin_5			(wallace_cout[59][5] ),
	.cin_6			(wallace_cout[59][6] ),
	.cin_7			(wallace_cout[59][7] ),
	.cin_8			(wallace_cout[59][8] ),
	.cin_9			(wallace_cout[59][9] ),
	.cin_10			(wallace_cout[59][10]),
	.cin_11			(wallace_cout[59][11]),
	.cin_12			(wallace_cout[59][12]),
	.cin_13			(wallace_cout[59][13]),
	.cin_14			(wallace_cout[59][14]),
	.cout_0			(wallace_cout[60][0] ),
	.cout_1			(wallace_cout[60][1] ),
	.cout_2			(wallace_cout[60][2] ),
	.cout_3			(wallace_cout[60][3] ),
	.cout_4			(wallace_cout[60][4] ),
	.cout_5			(wallace_cout[60][5] ),
	.cout_6			(wallace_cout[60][6] ),
	.cout_7			(wallace_cout[60][7] ),
	.cout_8			(wallace_cout[60][8] ),
	.cout_9			(wallace_cout[60][9] ),
	.cout_10		(wallace_cout[60][10]),
	.cout_11		(wallace_cout[60][11]),
	.cout_12		(wallace_cout[60][12]),
	.cout_13		(wallace_cout[60][13]),
	.cout_14		(wallace_cout[60][14]),
	.wallace_c		(wallace_c[60]       ),
	.wallace_s		(wallace_s[60]       )
);
wallace_tree wallace_tree_61(
	.wallace_input	(wallace_input[61]   ),
	.cin_0			(wallace_cout[60][0] ),
	.cin_1			(wallace_cout[60][1] ),
	.cin_2			(wallace_cout[60][2] ),
	.cin_3			(wallace_cout[60][3] ),
	.cin_4			(wallace_cout[60][4] ),
	.cin_5			(wallace_cout[60][5] ),
	.cin_6			(wallace_cout[60][6] ),
	.cin_7			(wallace_cout[60][7] ),
	.cin_8			(wallace_cout[60][8] ),
	.cin_9			(wallace_cout[60][9] ),
	.cin_10			(wallace_cout[60][10]),
	.cin_11			(wallace_cout[60][11]),
	.cin_12			(wallace_cout[60][12]),
	.cin_13			(wallace_cout[60][13]),
	.cin_14			(wallace_cout[60][14]),
	.cout_0			(wallace_cout[61][0] ),
	.cout_1			(wallace_cout[61][1] ),
	.cout_2			(wallace_cout[61][2] ),
	.cout_3			(wallace_cout[61][3] ),
	.cout_4			(wallace_cout[61][4] ),
	.cout_5			(wallace_cout[61][5] ),
	.cout_6			(wallace_cout[61][6] ),
	.cout_7			(wallace_cout[61][7] ),
	.cout_8			(wallace_cout[61][8] ),
	.cout_9			(wallace_cout[61][9] ),
	.cout_10		(wallace_cout[61][10]),
	.cout_11		(wallace_cout[61][11]),
	.cout_12		(wallace_cout[61][12]),
	.cout_13		(wallace_cout[61][13]),
	.cout_14		(wallace_cout[61][14]),
	.wallace_c		(wallace_c[61]       ),
	.wallace_s		(wallace_s[61]       )
);
wallace_tree wallace_tree_62(
	.wallace_input	(wallace_input[62]   ),
	.cin_0			(wallace_cout[61][0] ),
	.cin_1			(wallace_cout[61][1] ),
	.cin_2			(wallace_cout[61][2] ),
	.cin_3			(wallace_cout[61][3] ),
	.cin_4			(wallace_cout[61][4] ),
	.cin_5			(wallace_cout[61][5] ),
	.cin_6			(wallace_cout[61][6] ),
	.cin_7			(wallace_cout[61][7] ),
	.cin_8			(wallace_cout[61][8] ),
	.cin_9			(wallace_cout[61][9] ),
	.cin_10			(wallace_cout[61][10]),
	.cin_11			(wallace_cout[61][11]),
	.cin_12			(wallace_cout[61][12]),
	.cin_13			(wallace_cout[61][13]),
	.cin_14			(wallace_cout[61][14]),
	.cout_0			(wallace_cout[62][0] ),
	.cout_1			(wallace_cout[62][1] ),
	.cout_2			(wallace_cout[62][2] ),
	.cout_3			(wallace_cout[62][3] ),
	.cout_4			(wallace_cout[62][4] ),
	.cout_5			(wallace_cout[62][5] ),
	.cout_6			(wallace_cout[62][6] ),
	.cout_7			(wallace_cout[62][7] ),
	.cout_8			(wallace_cout[62][8] ),
	.cout_9			(wallace_cout[62][9] ),
	.cout_10		(wallace_cout[62][10]),
	.cout_11		(wallace_cout[62][11]),
	.cout_12		(wallace_cout[62][12]),
	.cout_13		(wallace_cout[62][13]),
	.cout_14		(wallace_cout[62][14]),
	.wallace_c		(wallace_c[62]       ),
	.wallace_s		(wallace_s[62]       )
);
wallace_tree wallace_tree_63(
	.wallace_input	(wallace_input[63]   ),
	.cin_0			(wallace_cout[62][0] ),
	.cin_1			(wallace_cout[62][1] ),
	.cin_2			(wallace_cout[62][2] ),
	.cin_3			(wallace_cout[62][3] ),
	.cin_4			(wallace_cout[62][4] ),
	.cin_5			(wallace_cout[62][5] ),
	.cin_6			(wallace_cout[62][6] ),
	.cin_7			(wallace_cout[62][7] ),
	.cin_8			(wallace_cout[62][8] ),
	.cin_9			(wallace_cout[62][9] ),
	.cin_10			(wallace_cout[62][10]),
	.cin_11			(wallace_cout[62][11]),
	.cin_12			(wallace_cout[62][12]),
	.cin_13			(wallace_cout[62][13]),
	.cin_14			(wallace_cout[62][14]),
	.cout_0			(wallace_cout[63][0] ),
	.cout_1			(wallace_cout[63][1] ),
	.cout_2			(wallace_cout[63][2] ),
	.cout_3			(wallace_cout[63][3] ),
	.cout_4			(wallace_cout[63][4] ),
	.cout_5			(wallace_cout[63][5] ),
	.cout_6			(wallace_cout[63][6] ),
	.cout_7			(wallace_cout[63][7] ),
	.cout_8			(wallace_cout[63][8] ),
	.cout_9			(wallace_cout[63][9] ),
	.cout_10		(wallace_cout[63][10]),
	.cout_11		(wallace_cout[63][11]),
	.cout_12		(wallace_cout[63][12]),
	.cout_13		(wallace_cout[63][13]),
	.cout_14		(wallace_cout[63][14]),
	.wallace_c		(wallace_c[63]       ),
	.wallace_s		(wallace_s[63]       )
);
wallace_tree wallace_tree_64(
	.wallace_input	(wallace_input[64]   ),
	.cin_0			(wallace_cout[63][0] ),
	.cin_1			(wallace_cout[63][1] ),
	.cin_2			(wallace_cout[63][2] ),
	.cin_3			(wallace_cout[63][3] ),
	.cin_4			(wallace_cout[63][4] ),
	.cin_5			(wallace_cout[63][5] ),
	.cin_6			(wallace_cout[63][6] ),
	.cin_7			(wallace_cout[63][7] ),
	.cin_8			(wallace_cout[63][8] ),
	.cin_9			(wallace_cout[63][9] ),
	.cin_10			(wallace_cout[63][10]),
	.cin_11			(wallace_cout[63][11]),
	.cin_12			(wallace_cout[63][12]),
	.cin_13			(wallace_cout[63][13]),
	.cin_14			(wallace_cout[63][14]),
	.cout_0			(wallace_cout[64][0] ),
	.cout_1			(wallace_cout[64][1] ),
	.cout_2			(wallace_cout[64][2] ),
	.cout_3			(wallace_cout[64][3] ),
	.cout_4			(wallace_cout[64][4] ),
	.cout_5			(wallace_cout[64][5] ),
	.cout_6			(wallace_cout[64][6] ),
	.cout_7			(wallace_cout[64][7] ),
	.cout_8			(wallace_cout[64][8] ),
	.cout_9			(wallace_cout[64][9] ),
	.cout_10		(wallace_cout[64][10]),
	.cout_11		(wallace_cout[64][11]),
	.cout_12		(wallace_cout[64][12]),
	.cout_13		(wallace_cout[64][13]),
	.cout_14		(wallace_cout[64][14]),
	.wallace_c		(wallace_c[64]       ),
	.wallace_s		(wallace_s[64]       )
);
wallace_tree wallace_tree_65(
	.wallace_input	(wallace_input[65]),
	.cin_0			(wallace_cout[64][0]),
	.cin_1			(wallace_cout[64][1]),
	.cin_2			(wallace_cout[64][2]),
	.cin_3			(wallace_cout[64][3]),
	.cin_4			(wallace_cout[64][4]),
	.cin_5			(wallace_cout[64][5]),
	.cin_6			(wallace_cout[64][6]),
	.cin_7			(wallace_cout[64][7]),
	.cin_8			(wallace_cout[64][8]),
	.cin_9			(wallace_cout[64][9]),
	.cin_10			(wallace_cout[64][10]),
	.cin_11			(wallace_cout[64][11]),
	.cin_12			(wallace_cout[64][12]),
	.cin_13			(wallace_cout[64][13]),
	.cin_14			(wallace_cout[64][14]),
	.cout_0			(),
	.cout_1			(),
	.cout_2			(),
	.cout_3			(),
	.cout_4			(),
	.cout_5			(),
	.cout_6			(),
	.cout_7			(),
	.cout_8			(),
	.cout_9			(),
	.cout_10		(),
	.cout_11		(),
	.cout_12		(),
	.cout_13		(),
	.cout_14		(),
	.wallace_c		(),
	.wallace_s		(wallace_s[65])
);

reg [65:0] add_c;
reg [65:0] add_s;
reg add_cin;
always @(posedge mul_clk)
begin
	if (~resetn) begin
		add_c <= 0;
		add_s <= 0;
		add_cin <= 0;
	end
	else begin
		add_c <= {wallace_c[64], wallace_c[63], wallace_c[62],
		          wallace_c[61], wallace_c[60], wallace_c[59],
		          wallace_c[58], wallace_c[57], wallace_c[56],
		          wallace_c[55], wallace_c[54], wallace_c[53],
		          wallace_c[52], wallace_c[51], wallace_c[50],
		          wallace_c[49], wallace_c[48], wallace_c[47],
		          wallace_c[46], wallace_c[45], wallace_c[44],
		          wallace_c[43], wallace_c[42], wallace_c[41],
		          wallace_c[40], wallace_c[39], wallace_c[38],
		          wallace_c[37], wallace_c[36], wallace_c[35],
		          wallace_c[34], wallace_c[33], wallace_c[32],
		          wallace_c[31], wallace_c[30], wallace_c[29],
		          wallace_c[28], wallace_c[27], wallace_c[26],
		          wallace_c[25], wallace_c[24], wallace_c[23],
		          wallace_c[22], wallace_c[21], wallace_c[20],
		          wallace_c[19], wallace_c[18], wallace_c[17],
		          wallace_c[16], wallace_c[15], wallace_c[14],
		          wallace_c[13], wallace_c[12], wallace_c[11],
		          wallace_c[10], wallace_c[9], wallace_c[8],
		          wallace_c[7], wallace_c[6], wallace_c[5],
		          wallace_c[4], wallace_c[3], wallace_c[2],
		          wallace_c[1], wallace_c[0], c[15]};
		add_s <= {wallace_s[65], wallace_s[64], wallace_s[63],
		          wallace_s[62], wallace_s[61], wallace_s[60],
		          wallace_s[59], wallace_s[58], wallace_s[57],
		          wallace_s[56], wallace_s[55], wallace_s[54],
		          wallace_s[53], wallace_s[52], wallace_s[51],
		          wallace_s[50], wallace_s[49], wallace_s[48],
		          wallace_s[47], wallace_s[46], wallace_s[45],
		          wallace_s[44], wallace_s[43], wallace_s[42],
		          wallace_s[41], wallace_s[40], wallace_s[39],
		          wallace_s[38], wallace_s[37], wallace_s[36],
		          wallace_s[35], wallace_s[34], wallace_s[33],
		          wallace_s[32], wallace_s[31], wallace_s[30],
		          wallace_s[29], wallace_s[28], wallace_s[27],
		          wallace_s[26], wallace_s[25], wallace_s[24],
		          wallace_s[23], wallace_s[22], wallace_s[21],
		          wallace_s[20], wallace_s[19], wallace_s[18],
		          wallace_s[17], wallace_s[16], wallace_s[15],
		          wallace_s[14], wallace_s[13], wallace_s[12],
		          wallace_s[11], wallace_s[10], wallace_s[9],
		          wallace_s[8], wallace_s[7], wallace_s[6],
		          wallace_s[5], wallace_s[4], wallace_s[3],
		          wallace_s[2], wallace_s[1], wallace_s[0]};
		add_cin <= c[16];
	end
end

wire [65:0] result_66bits;
assign result_66bits = add_c + add_s + add_cin;

assign result = result_66bits[63:0];
							
endmodule

module booth(
  input [65:0] x,
  input y0,
  input y1,
  input y2,
  output [65:0] p,
  output c
);
wire s_plus_2x;
wire s_minus_2x;
wire s_plus_x;
wire s_minus_x;
assign s_plus_2x = y0 & y1 & ~y2;
assign s_minus_2x = ~y0 & ~y1 & y2;
assign s_plus_x = y0 & ~y1 & ~y2 | ~y0 & y1 & ~y2;
assign s_minus_x = y0 & ~y1 & y2 | ~y0 & y1 & y2;

assign c = s_minus_x | s_minus_2x;
assign p = x & {66{s_plus_x}} | {x[64:0], 1'b0} & {66{s_plus_2x}}
         | ~x & {66{s_minus_x}} | {~x[64:0], 1'b1} & {66{s_minus_2x}};

endmodule

module wallace_tree(
	input [16:0] wallace_input,
	input cin_0,
	input cin_1,
	input cin_2,
	input cin_3,
	input cin_4,
	input cin_5,
	input cin_6,
	input cin_7,
	input cin_8,
	input cin_9,
	input cin_10,
	input cin_11,
	input cin_12,
	input cin_13,
	input cin_14,
	output cout_0,
	output cout_1,
	output cout_2,
	output cout_3,
	output cout_4,
	output cout_5,
	output cout_6,
	output cout_7,
	output cout_8,
	output cout_9,
	output cout_10,
	output cout_11,
	output cout_12,
	output cout_13,
	output cout_14,
	output wallace_c,
	output wallace_s
);
wire s_1_1;
wire s_1_2;
wire s_1_3;
wire s_1_4;
wire s_1_5;
wire s_1_6;
full_adder full_adder_1_1(
	.a		(wallace_input[0]	),
	.b		(wallace_input[1]	),
	.cin	(wallace_input[2]	),
	.cout	(cout_0				),
	.s		(s_1_1				)
);
full_adder full_adder_1_2(
	.a		(wallace_input[3]	),
	.b		(wallace_input[4]	),
	.cin	(wallace_input[5]	),
	.cout	(cout_1				),
	.s		(s_1_2				)
);
full_adder full_adder_1_3(
	.a		(wallace_input[6]	),
	.b		(wallace_input[7]	),
	.cin	(wallace_input[8]	),
	.cout	(cout_2				),
	.s		(s_1_3				)
);
full_adder full_adder_1_4(
	.a		(wallace_input[9]	),
	.b		(wallace_input[10]	),
	.cin	(wallace_input[11]	),
	.cout	(cout_3				),
	.s		(s_1_4				)
);
full_adder full_adder_1_5(
	.a		(wallace_input[12]	),
	.b		(wallace_input[13]	),
	.cin	(wallace_input[14]	),
	.cout	(cout_4				),
	.s		(s_1_5				)
);
half_adder half_adder_1_6(
	.a		(wallace_input[15]	),
	.b		(wallace_input[16]	),
	.cout	(cout_5				),
	.s		(s_1_6				)
);

wire s_2_1;
wire s_2_2;
wire s_2_3;
wire s_2_4;
full_adder full_adder_2_1(
	.a		(s_1_1				),
	.b		(s_1_2				),
	.cin	(s_1_3				),
	.cout	(cout_6				),
	.s		(s_2_1				)
);
full_adder full_adder_2_2(
	.a		(s_1_4				),
	.b		(s_1_5				),
	.cin	(s_1_6				),
	.cout	(cout_7				),
	.s		(s_2_2				)
);
full_adder full_adder_2_3(
	.a		(cin_0				),
	.b		(cin_1				),
	.cin	(cin_2				),
	.cout	(cout_8			),
	.s		(s_2_3				)
);
full_adder full_adder_2_4(
	.a		(cin_3				),
	.b		(cin_4				),
	.cin	(cin_5				),
	.cout	(cout_9				),
	.s		(s_2_4				)
);

wire s_3_1;
wire s_3_2;
full_adder full_adder_3_1(
	.a		(s_2_1				),
	.b		(s_2_2				),
	.cin	(s_2_3				),
	.cout	(cout_10			),
	.s		(s_3_1				)
);
full_adder full_adder_3_2(
	.a		(s_2_4				),
	.b		(cin_6				),
	.cin	(cin_7				),
	.cout	(cout_11			),
	.s		(s_3_2				)
);

wire s_4_1;
wire s_4_2;
full_adder full_adder_4_1(
	.a		(s_3_1				),
	.b		(s_3_2				),
	.cin	(cin_8				),
	.cout	(cout_12			),
	.s		(s_4_1				)
);
full_adder full_adder_4_2(
	.a		(cin_9				),
	.b		(cin_10				),
	.cin	(cin_11				),
	.cout	(cout_13			),
	.s		(s_4_2				)
);

wire s_5_1;
full_adder full_adder_5_1(
	.a		(s_4_1				),
	.b		(s_4_2				),
	.cin	(cin_12			),
	.cout	(cout_14			),
	.s		(s_5_1				)
);

full_adder full_adder_6_1(
	.a		(s_5_1				),
	.b		(cin_13			),
	.cin	(cin_14			),
	.cout	(wallace_c			),
	.s		(wallace_s			)
);

endmodule

module full_adder(
	input a,
	input b,
	input cin,
	output cout,
	output s
);
assign cout = b & cin | a & cin | a & b;
assign s = ~a & ~b & cin | ~a & b & ~cin | a & ~b & ~cin | a & b & cin;

endmodule

module half_adder(
	input a,
	input b,
	output cout,
	output s
);
assign cout = a & b;
assign s = ~a & b | a & ~b;

endmodule
